* NGSPICE file created from serv_0.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_1 D SE SI CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_ip_sram__sram256x8m8wm1 abstract view
.subckt gf180mcu_fd_ip_sram__sram256x8m8wm1 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7]
+ CEN CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] GWEN Q[0] Q[1] Q[2] Q[3] Q[4] Q[5]
+ Q[6] Q[7] WEN[0] WEN[1] WEN[2] WEN[3] WEN[4] WEN[5] WEN[6] WEN[7] VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

.subckt serv_0 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb[0] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] vdd vss
XFILLER_95_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2106_ _0354_ _0458_ _0448_ _0367_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2037_ _0392_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[45\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _2939_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2006__I0 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2084__B _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1996__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1748__A2 _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[34\] u_arbiter.i_wb_cpu_rdt\[31\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ u_scanchain_local.clk u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_64_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1920__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2259__B _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[68\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1436__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1739__A2 _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2724_ _0113_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2655_ _0044_ io_in[4] u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1606_ _1029_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2164__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2586_ _0822_ _0873_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1537_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _0926_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1468_ u_arbiter.i_wb_cpu_dbus_adr\[13\] _0926_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1399_ u_cpu.cpu.csr_imm _0851_ _0876_ u_cpu.cpu.immdec.imm24_20\[0\] _0888_ _0889_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_76_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1902__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2672__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1418__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1969__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2091__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[2\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2440_ _0728_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_97_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2146__A2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2371_ u_arbiter.i_wb_cpu_dbus_adr\[11\] u_arbiter.i_wb_cpu_dbus_adr\[12\] _0678_
+ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1409__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2082__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _0096_ io_in[4] u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2137__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2638_ _0002_ io_in[4] u_cpu.rf_ram_if.rdata0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2569_ u_arbiter.i_wb_cpu_rdt\[28\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _0799_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1896__B2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1896__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2695__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1820__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1757__I _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2128__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1887__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1639__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2300__A2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1940_ u_arbiter.i_wb_cpu_dbus_dat\[22\] _0286_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2064__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1871_ _0260_ _0262_ _1204_ _0263_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1662__I1 u_cpu.rf_ram.data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1811__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2423_ _1163_ _0713_ _0717_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1616__B u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2354_ _0679_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2285_ _0379_ _0433_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2166__C _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2055__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1802__A1 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1577__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1869__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2294__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1688__S _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2710__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2046__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2046__B2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2521__A2 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2070_ u_arbiter.i_wb_cpu_rdt\[5\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _0899_
+ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2285__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2972_ _2972_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ u_arbiter.i_wb_cpu_dbus_dat\[16\] _0286_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2588__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1854_ _0891_ _0221_ _0248_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1785_ _0897_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2406_ _0705_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2337_ _0858_ u_cpu.cpu.immdec.imm24_20\[0\] _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2268_ _1029_ _0605_ _1192_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2199_ _0535_ _0540_ _0543_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2733__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2028__B2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2028__A1 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2579__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2200__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2503__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[64\] u_scanchain_local.module_data_in\[63\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[26\] u_scanchain_local.clk u_scanchain_local.module_data_in\[64\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _1003_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2756__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2122_ _0397_ _0426_ _0401_ _0465_ _0379_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_6_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2053_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_74_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2217__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2955_ _2955_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2886_ _2886_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1906_ _0290_ _0291_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1837_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _0228_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1768_ _1078_ _1076_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1941__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1699_ _1132_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2249__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2127__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2629__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1932__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2779__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1463__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2740_ _0129_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2412__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2671_ _0060_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1622_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\] _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_126_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1553_ u_cpu.rf_ram_if.rcnt\[0\] _0849_ _0850_ u_cpu.rf_ram_if.wen0_r _1008_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_67_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1484_ u_arbiter.i_wb_cpu_dbus_adr\[17\] _0904_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2191__A3 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2105_ _0385_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2036_ _0367_ _0394_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1454__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2938_ _2938_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2869_ _2869_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_11_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2084__C _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[27\] u_arbiter.i_wb_cpu_rdt\[24\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1905__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2723_ _0112_ io_in[4] u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ _0043_ io_in[4] u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2585_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1605_ _0861_ _1056_ _1057_ _0855_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1536_ _0894_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1372__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1467_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _0937_ _0942_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1398_ _0886_ _0887_ _0851_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2185__B _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2019_ _0362_ _0379_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2624__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2405__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[23\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[38\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2817__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2615__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2091__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[35\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ _0687_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1409__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2606__A1 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2082__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2706_ _0095_ io_in[4] u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2637_ _0001_ io_in[4] u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2568_ _0811_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1519_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1896__A2 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2499_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _0718_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1974__S _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[58\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1584__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1639__A2 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1870_ u_arbiter.i_wb_cpu_dbus_dat\[1\] _0254_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1811__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2422_ _0713_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2353_ u_arbiter.i_wb_cpu_dbus_adr\[2\] u_arbiter.i_wb_cpu_dbus_adr\[3\] _0678_ _0679_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2127__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2284_ _0338_ _0479_ _0617_ _0369_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2055__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1999_ u_arbiter.i_wb_cpu_rdt\[15\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _0898_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2212__C1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2662__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1566__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[1\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2046__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2506__B1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2357__I0 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2285__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2971_ _2971_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2283__B _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ _0300_ _0301_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2685__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1796__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1853_ u_cpu.cpu.state.init_done _0228_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1784_ _1163_ _1188_ _1031_ u_arbiter.i_wb_cpu_dbus_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2596__I0 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1548__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ u_arbiter.i_wb_cpu_dbus_adr\[28\] u_arbiter.i_wb_cpu_dbus_adr\[29\] _1073_
+ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2336_ _0335_ _0624_ _0662_ _0369_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2267_ _1020_ _1077_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2198_ u_cpu.cpu.immdec.imm30_25\[0\] _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2276__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2028__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1787__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1539__A1 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2267__A2 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1490__A3 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2019__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1778__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2323__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[57\] u_scanchain_local.module_data_in\[56\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[19\] u_scanchain_local.clk u_scanchain_local.module_data_in\[57\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_67_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ _0355_ _0393_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2052_ _1189_ u_arbiter.i_wb_cpu_rdt\[11\] _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2954_ _2954_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2885_ _2885_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1905_ u_arbiter.i_wb_cpu_rdt\[8\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1836_ _0234_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2569__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1767_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _1070_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2194__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1941__A1 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1698_ u_cpu.rf_ram_if.rdata1\[2\] _1131_ _1010_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2700__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2319_ _0381_ _0646_ _0650_ _0382_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2850__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2249__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2185__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1932__A1 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2488__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[2\] u_arbiter.i_wb_cpu_ack io_in[3] u_arbiter.i_wb_cpu_dbus_sel\[0\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2412__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2670_ _0059_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1621_ _0852_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2176__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2723__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1923__A1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1552_ _0999_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1483_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] u_cpu.cpu.ctrl.o_ibus_adr\[16\] _0949_ _0954_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_28_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2104_ _0397_ _0387_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2035_ _0333_ _0381_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2100__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2937_ _2937_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2868_ _2868_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2190__C _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2799_ _0184_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2167__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1819_ u_cpu.cpu.state.o_cnt_r\[3\] u_cpu.cpu.state.o_cnt\[2\] _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[9\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2746__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1905__A1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1905__B2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2330__A1 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2291__B _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2722_ _0111_ io_in[4] u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2653_ _0042_ io_in[4] u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2149__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2584_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1604_ u_cpu.cpu.branch_op _1016_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1535_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] u_cpu.cpu.ctrl.o_ibus_adr\[29\] _0989_ _0993_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1635__B u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1466_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _0937_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _0941_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1397_ _0865_ _0868_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2018_ _0345_ _0368_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2185__C _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2769__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2312__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1455__B _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2303__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _0094_ io_in[4] u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2636_ _0000_ io_in[4] u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2567_ u_arbiter.i_wb_cpu_rdt\[27\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _0799_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2542__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1518_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] u_cpu.cpu.ctrl.o_ibus_adr\[24\] u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _0971_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_59_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2498_ _0756_ _0759_ _0760_ _1036_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1449_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _0925_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__B _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2058__B1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1820__A3 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2524__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2421_ _0711_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2352_ _1073_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2283_ _0352_ _0376_ _0616_ _0479_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2127__I1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[22\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[37\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2460__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2807__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1998_ _1189_ u_arbiter.i_wb_cpu_rdt\[14\] _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2212__C2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2619_ _0844_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_u_scanchain_local.scan_flop\[25\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2506__B2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2506__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2970_ _2970_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2283__C _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1921_ u_arbiter.i_wb_cpu_rdt\[14\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1852_ _0247_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1783_ _0852_ _1163_ _1031_ u_arbiter.i_wb_cpu_dbus_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1548__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2404_ _0704_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2335_ _1192_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2266_ _0856_ u_cpu.cpu.decode.opcode\[1\] _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2197_ _1192_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[48\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2433__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1787__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1490__A4 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__A2 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2120_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2051_ _0899_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_48_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2652__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2953_ _2953_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_90_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1904_ u_arbiter.i_wb_cpu_dbus_dat\[9\] _0286_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1769__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2884_ _2884_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1835_ _0892_ u_cpu.cpu.state.o_cnt_r\[2\] _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1766_ _1171_ _1177_ _1064_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_u_scanchain_local.scan_flop\[0\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1926__C1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1941__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1697_ _1128_ _0019_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2188__C _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2318_ _0381_ _0648_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2249_ _0339_ _0340_ _0343_ _0363_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2009__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1932__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2675__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2098__C _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1448__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1923__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1972__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1551_ u_cpu.rf_ram.data\[0\] _0999_ _1000_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1482_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _0949_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _0953_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2103_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_rdt\[5\] _0900_ _0456_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2034_ _0388_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ _2936_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2867_ _2867_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1818_ u_cpu.cpu.state.o_cnt_r\[3\] u_cpu.cpu.state.o_cnt\[2\] _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ _0183_ io_in[4] u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2167__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1882__I _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1749_ u_cpu.cpu.bufreg.lsb\[1\] _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2698__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1602__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1993__S _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1905__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1381__A3 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2094__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1841__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2721_ _0110_ io_in[4] u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2149__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2652_ _0041_ io_in[4] u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2583_ _0816_ _0818_ _0820_ _0872_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2840__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1603_ _0860_ _0853_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1534_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _0989_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _0992_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1465_ _0907_ _0939_ _0940_ u_arbiter.o_wb_cpu_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1396_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.genblk1.misalign_trap_sync_r
+ _0871_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2321__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2017_ _0367_ _0347_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2085__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1832__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2919_ _2919_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_91_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1596__B1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2312__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2076__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2713__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1823__A1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1674__I1 u_cpu.rf_ram.data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[32\] u_arbiter.i_wb_cpu_rdt\[29\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_64_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2000__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2303__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1471__B _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ _0093_ io_in[4] u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2635_ _0012_ io_in[4] u_cpu.rf_ram_if.rdata1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2566_ _0810_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1517_ _0907_ _0978_ _0979_ u_arbiter.o_wb_cpu_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1750__B1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2497_ _0756_ _1091_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1448_ _0905_ _0924_ _0925_ _0927_ u_arbiter.o_wb_cpu_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2736__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[6\]_SI u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1379_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2058__B2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2058__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2230__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1584__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1639__A4 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2049__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2342__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2221__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2420_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _1181_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2759__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2524__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2351_ _0677_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2282_ _0343_ _0388_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2288__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2460__B2 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1997_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1646__S0 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2618_ _0892_ u_cpu.rf_ram_if.rreq_r _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2549_ u_arbiter.i_wb_cpu_rdt\[18\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _0799_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2279__A1 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2203__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2506__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1493__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1920_ u_arbiter.i_wb_cpu_dbus_dat\[15\] _0286_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1851_ u_cpu.cpu.mem_bytecnt\[1\] _1075_ _0039_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1782_ u_cpu.cpu.bufreg.lsb\[1\] _1188_ _1031_ u_arbiter.i_wb_cpu_dbus_sel\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2403_ u_arbiter.i_wb_cpu_dbus_adr\[27\] u_arbiter.i_wb_cpu_dbus_adr\[28\] _1073_
+ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2334_ _0900_ u_arbiter.i_wb_cpu_rdt\[19\] _0381_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2265_ _0601_ _0602_ _0603_ _1165_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2196_ _1016_ _0536_ _1165_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1484__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[21\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1935__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[36\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2050_ _0362_ _0371_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1466__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2952_ _2952_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2415__B2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1903_ _0289_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2883_ _2883_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1834_ _0891_ _1102_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2179__B1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[20\]_D u_arbiter.i_wb_cpu_rdt\[17\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_1765_ _1173_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1926__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1696_ _1130_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[15\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2317_ _0337_ _0385_ _0401_ _0646_ _0379_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2248_ _0580_ _0581_ _0587_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2179_ u_cpu.cpu.immdec.imm24_20\[4\] _0498_ _0519_ _0405_ _0524_ _0525_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[22\]_SI u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[11\]_D u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1393__A1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1564__B u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2826__D _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[62\] u_scanchain_local.module_data_in\[61\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[24\] u_scanchain_local.clk u_scanchain_local.module_data_in\[62\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA_u_scanchain_local.scan_flop\[9\]_D u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2350__S _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1550_ u_arbiter.i_wb_cpu_dbus_we _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[38\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1384__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1481_ _0952_ u_arbiter.o_wb_cpu_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2102_ _0863_ _0407_ _0455_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2033_ _0360_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1649__B _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2935_ _2935_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2866_ _2866_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1817_ _0222_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2797_ _0182_ io_in[4] u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1748_ _0878_ _0026_ _1160_ u_cpu.rf_ram.addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1679_ _1120_ u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1403__I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1602__A2 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2642__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2792__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2409__I u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2618__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1841__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2720_ _0109_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2651_ _0040_ io_in[4] u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1602_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.genblk1.misalign_trap_sync_r
+ _0857_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_2582_ _0858_ u_arbiter.i_wb_cpu_dbus_we u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _0869_
+ _0818_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1533_ _0907_ _0990_ _0991_ u_arbiter.o_wb_cpu_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1372__A4 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1464_ u_arbiter.i_wb_cpu_dbus_adr\[12\] _0905_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1395_ u_cpu.cpu.immdec.imm19_12_20\[6\] _0851_ _0876_ u_cpu.cpu.immdec.imm24_20\[2\]
+ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2609__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2016_ _0376_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2085__A2 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1832__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2918_ _2918_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2665__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1596__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2849_ u_cpu.rf_ram_if.wdata1_r\[2\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1899__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1842__B _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2076__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1823__A2 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1587__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2000__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[25\] u_arbiter.i_wb_cpu_rdt\[22\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2303__A3 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2688__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2703_ _0092_ io_in[4] u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2634_ _0011_ io_in[4] u_cpu.rf_ram_if.rdata1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2565_ u_arbiter.i_wb_cpu_rdt\[26\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _0799_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1516_ u_arbiter.i_wb_cpu_dbus_adr\[25\] _0926_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2496_ u_cpu.cpu.ctrl.i_jump _1081_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1750__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1447_ u_arbiter.i_wb_cpu_dbus_adr\[8\] _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1378_ _0863_ _0865_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2058__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1569__A1 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A3 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1999__S _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2297__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2049__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2830__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2509__B1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2524__A3 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2350_ u_cpu.cpu.alu.cmp_r _0244_ _1029_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2281_ u_cpu.cpu.csr_imm _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2288__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1799__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2460__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1996_ _0350_ _0352_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1646__S1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1971__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2617_ _0851_ _0843_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2703__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2548_ _0801_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2479_ _0748_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_29_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2853__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2279__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2451__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2203__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ _0237_ _0246_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2353__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1781_ u_cpu.cpu.bne_or_bge _0852_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2726__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2402_ _0703_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2333_ _0900_ _0272_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2264_ u_cpu.cpu.immdec.imm7 _0407_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2195_ u_cpu.cpu.immdec.imm30_25\[1\] _0407_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2130__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2433__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2197__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1979_ _0339_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2121__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2424__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2749__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2173__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2188__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1935__A1 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2951_ _2951_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1902_ u_arbiter.i_wb_cpu_rdt\[7\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[8\] _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2882_ _2882_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1833_ _0233_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2179__B2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2179__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1926__A1 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1764_ _0856_ _1022_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1926__B2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1695_ u_cpu.rf_ram_if.rdata1\[1\] _1129_ _1010_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2316_ _0337_ _0626_ _0647_ _0621_ _0402_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ u_cpu.cpu.immdec.imm7 _1170_ _0544_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2178_ _0498_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1614__B1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1393__A2 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[55\] u_scanchain_local.module_data_in\[54\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[17\] u_scanchain_local.clk u_scanchain_local.module_data_in\[55\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1384__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1480_ u_arbiter.i_wb_cpu_dbus_adr\[16\] _0951_ _0894_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2333__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2101_ _0405_ _0446_ _0450_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2032_ _1189_ u_arbiter.i_wb_cpu_rdt\[15\] _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1710__S _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2934_ _2934_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1649__C _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2865_ _2865_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_11_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1816_ _0891_ _0221_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2021__B1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2796_ _0181_ io_in[4] u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1375__A2 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1747_ _0879_ _1001_ _1158_ _1162_ u_cpu.rf_ram.addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1678_ u_cpu.rf_ram_if.wdata0_r\[1\] u_cpu.rf_ram_if.wdata1_r\[1\] _0998_ _1120_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2324__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[20\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2088__B1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[35\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1602__A3 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2260__B1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2315__A1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[0\] io_in[2] io_in[3] u_arbiter.o_wb_cpu_cyc u_scanchain_local.clk
+ u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_92_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2650_ _0039_ io_in[4] u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2361__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1601_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.init_done _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2581_ _0819_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1532_ u_arbiter.i_wb_cpu_dbus_adr\[29\] _0926_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1463_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _0937_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2306__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1394_ u_cpu.cpu.immdec.imm19_12_20\[5\] u_cpu.rf_ram_if.rtrig0 _0883_ _0884_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2015_ _0360_ _0371_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2490__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2917_ _2917_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_52_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2848_ u_cpu.rf_ram_if.wdata1_r\[1\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2779_ _0165_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1414__I _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1520__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[28\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2536__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[18\] u_arbiter.i_wb_cpu_rdt\[15\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_75_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2472__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ _0091_ io_in[4] u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2633_ _0010_ io_in[4] u_cpu.rf_ram_if.rdata1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2564_ _0809_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2527__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1515_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2495_ u_cpu.cpu.ctrl.i_jump _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1750__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1446_ _0904_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1377_ _0859_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1502__A2 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2632__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2782__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1569__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2509__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2509__B2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1763__B _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2280_ _0613_ _0607_ _0614_ _0445_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2655__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2445__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1995_ _0354_ _0355_ _0356_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_140_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1420__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1971__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2616_ _1011_ _0843_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2547_ u_arbiter.i_wb_cpu_rdt\[17\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _0799_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2478_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[25\]
+ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1429_ _0907_ _0911_ _0912_ u_arbiter.o_wb_cpu_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2678__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1478__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1780_ _0886_ _1187_ _1165_ u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2589__B _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2401_ u_arbiter.i_wb_cpu_dbus_adr\[26\] u_arbiter.i_wb_cpu_dbus_adr\[27\] _1073_
+ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2332_ _0411_ _0479_ _0449_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1713__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2263_ _1165_ _0584_ _0382_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2194_ _0333_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1469__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2130__A2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1641__A1 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1978_ u_arbiter.i_wb_cpu_rdt\[8\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _0899_
+ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2820__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1422__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2121__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2188__A2 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1935__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2428__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2112__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ _2950_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2881_ _2881_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1901_ _0287_ _0288_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1623__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1832_ _0892_ u_cpu.cpu.state.o_cnt_r\[0\] _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2843__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2179__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1763_ _1174_ _1068_ _1091_ _0857_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1926__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1694_ _1128_ _0018_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2112__B _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2315_ _0449_ _0479_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2246_ _0582_ _0583_ _0585_ _1170_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2177_ u_cpu.cpu.immdec.imm30_25\[0\] _0333_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1862__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[61\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1398__B _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1614__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1917__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2590__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2716__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1853__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1605__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[48\] u_scanchain_local.module_data_in\[47\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[10\] u_scanchain_local.clk u_scanchain_local.module_data_in\[48\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2030__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2333__A2 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2359__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _0333_ _0403_ _0452_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_2031_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2097__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2933_ _2933_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2864_ _2864_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2795_ _0180_ io_in[4] u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1815_ _1014_ _1195_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2021__A1 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2021__B2 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1746_ u_cpu.cpu.immdec.imm11_7\[4\] _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1677_ _1119_ u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2739__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2324__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2229_ _0479_ _0481_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2088__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1835__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1686__I1 u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2260__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2260__B2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2012__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2315__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2079__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1826__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2251__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1766__B _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ _0852_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ _0817_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1531_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1462_ _0905_ _0935_ _0937_ _0938_ u_arbiter.o_wb_cpu_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_84_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2306__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1393_ u_cpu.rf_ram_if.rtrig0 _0862_ _0881_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_80_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1721__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2014_ _0372_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1668__I1 u_cpu.rf_ram.data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2490__B2 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2916_ _2916_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_91_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2847_ _0214_ io_in[4] u_cpu.rf_ram_if.rcnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2778_ _0164_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1729_ u_cpu.raddr\[0\] _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2300__B _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1587__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2536__A2 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2701_ _0090_ io_in[4] u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _0009_ io_in[4] u_cpu.rf_ram_if.rdata1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2563_ u_arbiter.i_wb_cpu_rdt\[25\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _0799_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1514_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] u_cpu.cpu.ctrl.o_ibus_adr\[23\] _0971_ _0977_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _1106_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[34\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1445_ _0922_ _0923_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1376_ _0854_ _0861_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1502__A3 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2547__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[49\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1569__A3 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2518__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[30\] u_arbiter.i_wb_cpu_rdt\[27\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1763__C _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2367__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1496__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ u_arbiter.i_wb_cpu_rdt\[2\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] _0898_
+ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1956__B1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1420__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2615_ _1128_ _0024_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[18\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2546_ _0800_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2477_ _0747_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1428_ u_arbiter.i_wb_cpu_dbus_adr\[4\] _0905_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1359_ u_cpu.rf_ram_if.rcnt\[0\] _0849_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[32\]_D u_arbiter.i_wb_cpu_rdt\[29\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1938__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0702_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2331_ _0607_ _0659_ _0660_ _0661_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2262_ _0338_ _0405_ _0600_ _0395_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2193_ _1029_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2772__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[23\]_D u_arbiter.i_wb_cpu_rdt\[20\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1929__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _0335_ _0336_ _0337_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_14_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2529_ _0402_ _0783_ _0787_ _0336_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_121_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[14\]_D u_arbiter.i_wb_cpu_rdt\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2645__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1396__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2795__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2880_ _2880_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1900_ u_arbiter.i_wb_cpu_rdt\[6\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1623__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _0229_ _0232_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1387__A1 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1762_ _1016_ u_cpu.cpu.decode.opcode\[1\] _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1693_ u_cpu.rf_ram.regzero _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2314_ u_arbiter.i_wb_cpu_rdt\[17\] u_arbiter.i_wb_cpu_rdt\[1\] _0899_ _0646_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2245_ _0584_ _0583_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2176_ _0395_ _0518_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2555__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1862__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1614__A2 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1378__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1853__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2405__I1 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1369__A1 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1541__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2030_ _0334_ _0389_ _0390_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2097__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2375__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1844__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2810__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2932_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2863_ _2863_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1719__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2794_ _0179_ io_in[4] u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1814_ _1207_ _0220_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1745_ _0877_ _1001_ _1161_ u_cpu.rf_ram.addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1676_ u_cpu.rf_ram_if.wdata0_r\[0\] u_cpu.rf_ram_if.wdata1_r\[0\] _0998_ _1119_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1780__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1532__A1 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2228_ _0336_ _0388_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2159_ _0470_ _0469_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2260__A2 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2012__A2 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1771__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2571__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2323__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2833__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1826__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[60\] u_scanchain_local.module_data_in\[59\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[22\] u_scanchain_local.clk u_scanchain_local.module_data_in\[60\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\] u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _0980_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1782__B _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1762__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1461_ u_arbiter.i_wb_cpu_dbus_adr\[11\] _0926_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1392_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _0859_ _0866_ _0882_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_45_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[51\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2314__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ _0339_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2490__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2915_ _2915_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2846_ u_cpu.rf_ram_if.rtrig0 io_in[4] u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2777_ _0163_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2706__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ _1001_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1753__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1659_ _0886_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1505__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2553__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2300__C _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2856__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1992__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1744__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2210__C _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2472__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2729__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _0089_ io_in[4] u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2631_ _0008_ io_in[4] u_cpu.rf_ram_if.rdata1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2562_ _0808_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1513_ _0907_ _0975_ _0976_ u_arbiter.o_wb_cpu_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1735__A1 u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2493_ _0873_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1444_ _0922_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2160__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1375_ _0864_ u_cpu.cpu.decode.op26 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2563__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ _0021_ io_in[4] u_cpu.rf_ram.rdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2518__A3 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[23\] u_arbiter.i_wb_cpu_rdt\[20\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2142__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2445__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2383__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1993_ u_arbiter.i_wb_cpu_rdt\[4\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] _0898_
+ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ _0719_ _0841_ _0842_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2545_ u_arbiter.i_wb_cpu_rdt\[16\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2476_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[24\]
+ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1427_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2133__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1358_ u_cpu.rf_ram_if.rcnt\[1\] _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2124__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2124__B2 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1478__A3 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[33\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1938__A1 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[48\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ u_cpu.cpu.immdec.imm19_12_20\[7\] _0607_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2261_ _0598_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2115__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2192_ _1016_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1976_ u_arbiter.i_wb_cpu_rdt\[7\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _0897_
+ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1929__A1 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2528_ _0368_ _0388_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2459_ _0718_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2106__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1865__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2036__B _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1632__A3 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1875__B _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1396__A2 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2593__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[2\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ _0892_ _1165_ _0231_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1761_ u_cpu.cpu.bufreg.c_r _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1387__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1692_ _1127_ u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2336__B2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2336__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2313_ _0607_ _0643_ _0644_ _0645_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2244_ u_cpu.cpu.immdec.imm31 _1020_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2175_ _0368_ _0350_ _0402_ _0520_ _0403_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_54_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2571__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1959_ u_arbiter.i_wb_cpu_rdt\[28\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[29\] _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_66_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2327__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1369__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2762__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2318__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2931_ _2931_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2391__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2862_ _2862_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_54_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2793_ _0178_ io_in[4] u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1813_ u_cpu.raddr\[1\] _0217_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1744_ u_cpu.cpu.immdec.imm11_7\[3\] _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1780__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1675_ _1118_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1532__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2227_ _0361_ _0567_ _0379_ _0385_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2158_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_rdt\[7\] _0899_ _0505_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2635__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2089_ _0360_ _0380_ _0443_ _0408_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2785__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1771__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2323__I1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[53\] u_scanchain_local.module_data_in\[52\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[15\] u_scanchain_local.clk u_scanchain_local.module_data_in\[53\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2539__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1762__A2 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1460_ _0929_ _0922_ _0923_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1391_ u_cpu.cpu.immdec.imm24_20\[1\] _0874_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2658__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2314__I1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2012_ _1189_ u_arbiter.i_wb_cpu_rdt\[8\] _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2914_ _2914_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_52_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2134__B _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2845_ _0213_ io_in[4] u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2776_ _0162_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1727_ u_cpu.rf_ram_if.rcnt\[0\] u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[2\]
+ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1658_ _1048_ _1095_ _1096_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1753__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1589_ _1041_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2466__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2309__B _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2069__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2218__B1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1441__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1992__A2 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2800__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2457__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2630_ _0007_ io_in[4] u_cpu.rf_ram_if.rdata1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2561_ u_arbiter.i_wb_cpu_rdt\[24\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _0799_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1512_ u_arbiter.i_wb_cpu_dbus_adr\[24\] _0926_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1735__A2 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2492_ _0864_ _0870_ _0866_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1443_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _0913_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1374_ u_cpu.cpu.decode.op21 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2129__B _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1959__C1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2828_ _0020_ io_in[4] u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2759_ _0145_ io_in[4] u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2823__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2439__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1878__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[41\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[16\] u_arbiter.i_wb_cpu_rdt\[13\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_93_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1653__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1992_ _0899_ _0272_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2846__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1405__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1956__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2412__B _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2613_ u_cpu.cpu.state.ibus_cyc _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2544_ _1190_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2475_ _0746_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1426_ _0900_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] u_cpu.cpu.ctrl.o_ibus_adr\[2\] _0910_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1357_ u_cpu.rf_ram_if.rcnt\[2\] _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_97_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[64\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2124__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2719__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1883__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1938__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2060__A1 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2260_ _0397_ _0356_ _0401_ _0338_ _0379_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2115__A2 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2191_ _0855_ _0857_ u_arbiter.i_wb_cpu_dbus_we _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_19_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ u_arbiter.i_wb_cpu_rdt\[9\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] _0897_
+ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1929__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2051__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2142__B _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2569__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2527_ u_cpu.cpu.immdec.imm11_7\[3\] _0763_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2458_ _0737_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_130_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1409_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0894_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2389_ u_arbiter.i_wb_cpu_dbus_adr\[20\] u_arbiter.i_wb_cpu_dbus_adr\[21\] _1073_
+ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1865__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1865__B2 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2290__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2042__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1396__A3 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[9\] u_arbiter.i_wb_cpu_rdt\[6\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_48_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1856__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2691__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1608__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2227__B _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2033__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1760_ u_cpu.cpu.alu.i_rs1 _1168_ _1170_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1691_ u_cpu.rf_ram_if.wdata1_r\[7\] u_cpu.cpu.o_wdata0 _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2389__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2336__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2312_ u_cpu.cpu.immdec.imm19_12_20\[5\] _0607_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2243_ _0855_ _1016_ u_cpu.cpu.decode.opcode\[1\] _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2174_ _0335_ _0397_ _0401_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1958_ _0324_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1889_ _1204_ _0252_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2327__A2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[32\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1838__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1730__I _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[47\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2263__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2015__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2930_ _2930_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2254__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2861_ _2861_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1812_ _0219_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2792_ _0177_ io_in[4] u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1743_ _1158_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1674_ u_cpu.rf_ram.rdata\[7\] u_cpu.rf_ram.data\[7\] _0026_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2190__B1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2226_ _1189_ u_arbiter.i_wb_cpu_rdt\[13\] _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1550__I u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2493__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2157_ _0503_ _0498_ _0504_ _0476_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2088_ _0355_ _0425_ _0409_ _0442_ _0438_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2236__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2539__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_scanchain_local.scan_flop\[46\] u_scanchain_local.module_data_in\[45\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[8\] u_scanchain_local.clk u_scanchain_local.module_data_in\[46\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1390_ _0877_ _0878_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2011_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2227__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2913_ _2913_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_52_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2134__C _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2844_ _0212_ io_in[4] u_cpu.rf_ram_if.rdata0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2775_ _0161_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1726_ _1148_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1657_ _0041_ _1101_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1588_ _1014_ u_cpu.cpu.genblk3.csr.mcause31 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1910__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2209_ _0354_ _0370_ _0347_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2752__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2218__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2218__B2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2325__B _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2060__B _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[2\]_D u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2209__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1432__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2560_ _0807_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2625__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1511_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2491_ _0754_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1735__A3 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1442_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2397__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2775__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1373_ u_cpu.cpu.decode.co_ebreak _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1959__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ _0019_ io_in[4] u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2758_ _0015_ io_in[4] u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1709_ _1128_ _0023_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2689_ _0078_ io_in[4] u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2611__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2648__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1973__I0 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2798__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1991_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _0382_ _0228_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2543_ _0891_ _0798_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2474_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1425_ _0907_ _0908_ _0909_ u_arbiter.o_wb_cpu_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_u_scanchain_local.scan_flop\[26\]_D u_arbiter.i_wb_cpu_rdt\[23\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1580__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1733__I _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1635__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[17\]_D u_arbiter.i_wb_cpu_rdt\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1399__A1 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1399__B2 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2060__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1571__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2190_ _0531_ _0533_ _0534_ _0381_ _0382_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1874__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2813__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1974_ u_arbiter.i_wb_cpu_rdt\[10\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _0897_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2051__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1562__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2526_ _1162_ _0763_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2457_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1408_ _0895_ u_arbiter.o_wb_cpu_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[31\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2388_ _0696_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1865__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3009_ io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2317__C _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2042__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1664__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1891__C _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2836__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2353__I0 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1856__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2508__B _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1608__A2 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2227__C _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2243__B u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1690_ _0998_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[54\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1373__I u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2311_ u_cpu.cpu.immdec.imm19_12_20\[6\] _1192_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2242_ u_cpu.cpu.immdec.imm19_12_20\[0\] _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2173_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_rdt\[8\] _0900_ _0519_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1957_ u_arbiter.i_wb_cpu_rdt\[27\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[28\] _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2709__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1888_ _1196_ _0277_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1783__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2509_ _0397_ _0354_ _0401_ _0340_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2015__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1774__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1829__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2254__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2860_ _2860_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_30_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1811_ _1193_ _1206_ _0217_ _0218_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_15_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1368__I _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2791_ _0013_ io_in[4] u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1742_ _0885_ _1001_ _1158_ _1159_ u_cpu.rf_ram.addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ _1117_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1517__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2565__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2190__B2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2225_ _0900_ u_arbiter.i_wb_cpu_rdt\[29\] _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2493__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2156_ u_cpu.cpu.immdec.imm24_20\[3\] _0496_ _0382_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2087_ _0350_ _0352_ _0414_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ _2989_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2681__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1756__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2103__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2236__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1995__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1747__B2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2547__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[39\] u_scanchain_local.module_data_in\[38\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[1\] u_scanchain_local.clk u_scanchain_local.module_data_in\[39\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_136_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2172__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2010_ _0370_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2912_ _2912_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_143_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1986__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2843_ _0211_ io_in[4] u_cpu.rf_ram_if.rdata1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[31\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2774_ _0160_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1725_ u_cpu.rf_ram_if.rdata0\[7\] _1139_ u_cpu.rf_ram_if.rtrig0 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1738__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[46\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2150__C _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1656_ _1106_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1587_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\]
+ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2163__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1910__A1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2466__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2208_ _0340_ _0393_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2139_ _0480_ _0488_ _0489_ _0345_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2218__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1672__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2154__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2457__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2209__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1968__A1 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1510_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _0971_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2490_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1441_ _0907_ _0920_ _0921_ u_arbiter.o_wb_cpu_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1372_ _0854_ u_cpu.cpu.decode.op21 _0859_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_64_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__A1 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2826_ _0018_ io_in[4] u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1556__I _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2757_ _0016_ io_in[4] u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2688_ _0077_ io_in[4] u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1708_ _1138_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1639_ _0860_ _0854_ u_cpu.cpu.alu.cmp_r _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_67_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2439__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1973__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[5\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1990_ _1189_ u_arbiter.i_wb_cpu_rdt\[5\] _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2611_ _0891_ u_cpu.cpu.genblk3.csr.timer_irq_r _0676_ _0840_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2742__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2542_ _0900_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2473_ _0745_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2118__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1424_ u_arbiter.i_wb_cpu_dbus_adr\[3\] _0905_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2156__B _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1487__S _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2809_ _0194_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2109__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1399__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2765__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[21\] u_arbiter.i_wb_cpu_rdt\[18\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_3_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2371__I1 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2520__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1973_ u_arbiter.i_wb_cpu_rdt\[11\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _0897_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2587__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2339__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2525_ _0764_ _0781_ _0782_ _0784_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2456_ _0736_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1562__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1407_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2387_ u_arbiter.i_wb_cpu_dbus_adr\[19\] u_arbiter.i_wb_cpu_dbus_adr\[20\] _1073_
+ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2511__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2638__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3008_ io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2788__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2578__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1680__S _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2502__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[69\] u_scanchain_local.module_data_in\[68\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[31\] u_scanchain_local.clk u_scanchain_local.module_data_in\[69\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2310_ _0381_ _0631_ _0642_ _0382_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_3_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2241_ u_cpu.cpu.immdec.imm30_25\[5\] _0542_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2172_ _0350_ _0416_ _0507_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2257__B1 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1956_ _0321_ _0282_ _0286_ _0322_ _0323_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2153__C _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1887_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _1197_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1783__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2508_ _0402_ _0768_ _0404_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2439_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[6\]
+ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2328__C _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2803__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2023__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2238__C _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1462__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1810_ u_cpu.raddr\[0\] _0216_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_15_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_scanchain_local.scan_flop\[21\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2790_ _0176_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1741_ u_cpu.cpu.immdec.imm11_7\[2\] _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1765__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1672_ u_cpu.rf_ram.rdata\[6\] u_cpu.rf_ram.data\[6\] _0026_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2478__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2224_ _0562_ _0564_ _0565_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2155_ u_cpu.cpu.immdec.imm24_20\[2\] _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2086_ _1031_ _0407_ _0441_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2164__B _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1453__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2988_ _2988_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2826__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1939_ _0311_ _0312_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1756__A2 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1508__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2181__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2058__C _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[44\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1995__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1747__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2249__B _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2911_ _2911_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_44_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2849__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_cpu.rf_ram.RAM0_A[7] u_cpu.rf_ram.addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1986__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1379__I u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2842_ u_cpu.rf_ram_if.wtrig0 io_in[4] u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2235__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2773_ _0159_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1724_ _1147_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1655_ _0857_ _1016_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1586_ u_cpu.cpu.state.o_cnt_r\[3\] _1037_ _1038_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2163__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1910__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2207_ _0340_ _0433_ _0549_ _0401_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[67\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2138_ _0356_ _0370_ _0393_ _0338_ _0347_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2069_ u_arbiter.i_wb_cpu_rdt\[6\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] _0899_
+ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1426__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1977__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1417__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1968__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2090__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2217__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[51\] u_scanchain_local.module_data_in\[50\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[13\] u_scanchain_local.clk u_scanchain_local.module_data_in\[51\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_51_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1440_ u_arbiter.i_wb_cpu_dbus_adr\[7\] _0905_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xu_scanchain_local.out_flop u_scanchain_local.module_data_in\[69\] u_scanchain_local.clk
+ u_scanchain_local.data_out_i vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__2145__A2 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1371_ _0860_ u_cpu.cpu.bne_or_bge _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2671__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1959__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2081__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2825_ _0017_ io_in[4] u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2756_ _0144_ io_in[4] u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2687_ _0076_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1707_ u_cpu.rf_ram_if.rdata1\[5\] _1137_ _1010_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1638_ u_cpu.cpu.state.o_cnt_r\[0\] _1038_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1569_ _1005_ _1012_ _1013_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_24_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1895__A1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2072__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1670__I1 u_cpu.rf_ram.data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1886__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2694__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[30\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1638__A1 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[45\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2063__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2610_ u_cpu.cpu.genblk3.csr.o_new_irq _0228_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2541_ u_arbiter.i_wb_cpu_ack u_arbiter.o_wb_cpu_adr\[1\] _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2472_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2118__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1423_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _0902_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1877__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1629__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2054__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1801__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2808_ _0193_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2739_ _0128_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2109__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1868__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2293__B2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2045__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1678__S _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__A2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[14\] u_arbiter.i_wb_cpu_rdt\[11\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1859__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2284__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2036__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2587__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2524_ _0407_ _0337_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2455_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[14\]
+ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1562__A3 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2386_ _0695_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1406_ _0893_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3007_ io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_43_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2027__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2732__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2266__A1 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2018__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2240_ _0405_ _0575_ _0579_ _1192_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2171_ _0335_ _0388_ _0367_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[7] u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2257__B2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2257__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1955_ u_arbiter.i_wb_cpu_rdt\[26\] _1204_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1886_ _0272_ _0273_ _0275_ _0276_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2507_ _0374_ _0593_ _0635_ _0767_ _0408_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2438_ _0727_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_29_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2755__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2369_ u_arbiter.i_wb_cpu_dbus_adr\[10\] u_arbiter.i_wb_cpu_dbus_adr\[11\] _0678_
+ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2420__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[7\] u_arbiter.i_wb_cpu_rdt\[4\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_43_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2628__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1740_ _1126_ _0886_ _1001_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1671_ _1116_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2270__B _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2175__B1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2778__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2223_ _0382_ _0404_ _0559_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2154_ _0464_ _0502_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2085_ _0371_ _0404_ _0440_ _1192_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_4_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2164__C _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ _2987_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1938_ u_arbiter.i_wb_cpu_rdt\[20\] _0273_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1869_ _0252_ _0261_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1913__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1686__S _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1995__A3 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[5\]_D u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1380__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2249__C _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2910_ _2910_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_91_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[6] u_cpu.rf_ram.addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2841_ u_cpu.cpu.o_wdata0 io_in[4] u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2235__I1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2772_ _0158_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1723_ u_cpu.rf_ram_if.rdata0\[6\] _1137_ u_cpu.rf_ram_if.rtrig0 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1994__I0 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1654_ _1104_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1585_ u_cpu.cpu.decode.op26 _0867_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1371__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2206_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_rdt\[11\] _0900_ _0549_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2137_ _0338_ _0388_ _0393_ _0427_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2068_ _0372_ _0375_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2623__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1977__A3 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1362__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[11\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2090__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2217__I1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[44\] u_scanchain_local.module_data_in\[43\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[6\] u_scanchain_local.clk u_scanchain_local.module_data_in\[44\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1370_ u_cpu.cpu.decode.co_mem_word _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2816__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[38\]_D u_scanchain_local.module_data_in\[37\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2081__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2824_ _0209_ io_in[4] u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2755_ _0143_ io_in[4] u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2686_ _0075_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1706_ _1128_ _0022_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1637_ _0853_ _1087_ _1088_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_63_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[34\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1568_ u_arbiter.i_wb_cpu_dbus_we _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1499_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1895__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1647__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1802__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[29\]_D u_arbiter.i_wb_cpu_rdt\[26\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2072__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2839__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1886__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1638__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2063__A2 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ _0580_ _0796_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[57\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2471_ _0744_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_5_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1422_ _0904_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2054__A2 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1801__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2807_ _0192_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2738_ _0127_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1565__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2669_ _0058_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1868__A2 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2293__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2045__A2 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2661__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1859__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2284__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1971_ u_arbiter.i_wb_cpu_ack _0894_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2273__B _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2036__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1795__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2587__A3 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2523_ _0470_ _0363_ _0404_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1547__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2454_ _0735_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_116_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2385_ u_arbiter.i_wb_cpu_dbus_adr\[18\] u_arbiter.i_wb_cpu_dbus_adr\[19\] _1073_
+ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1405_ _0892_ u_cpu.cpu.state.ibus_cyc _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_25_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2167__C _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3006_ _3006_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2027__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1578__I u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1786__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2684__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2403__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_scanchain_local.scan_flop\[44\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[59\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2266__A2 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2018__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1777__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1529__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2268__B _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ _0498_ _0514_ _0515_ _0516_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_59_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[6] u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2257__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1954_ u_arbiter.i_wb_cpu_dbus_dat\[27\] _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1885_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _0268_ _0257_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2193__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ _0340_ _0370_ _0393_ _0354_ _0593_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2437_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2368_ _0686_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2299_ _0401_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1759__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2420__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2559__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1998__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1462__A3 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2411__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1670_ u_cpu.rf_ram.rdata\[5\] u_cpu.rf_ram.data\[5\] _0026_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2175__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2478__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2222_ u_cpu.cpu.immdec.imm30_25\[3\] _0539_ _0563_ u_cpu.cpu.immdec.imm30_25\[4\]
+ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2153_ u_cpu.cpu.immdec.imm24_20\[2\] _0496_ _0501_ _0334_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2084_ _0408_ _0439_ _0399_ _0404_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1989__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2986_ _2986_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1937_ u_arbiter.i_wb_cpu_dbus_dat\[21\] _0286_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1868_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[1\] _1196_ _0261_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1799_ _1196_ _1199_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2166__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2722__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1913__A1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2157__B2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1380__A2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[8\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[5] u_cpu.rf_ram.addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1691__I0 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2840_ u_cpu.rf_ram_if.wdata0_r\[6\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1435__A3 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2771_ _0157_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2745__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1722_ _1146_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1609__C u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1653_ u_arbiter.i_wb_cpu_ibus_adr\[0\] u_cpu.cpu.ctrl.pc_plus_4_cy_r _1105_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1584_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\]
+ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_63_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1371__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2205_ _0526_ _0546_ _0547_ _0530_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2320__A1 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2136_ _0484_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2067_ u_cpu.cpu.bne_or_bge _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__A4 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2969_ _2969_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2139__B2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1362__A2 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2085__C _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2768__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[37\] u_scanchain_local.module_data_in\[36\] io_in[3]
+ u_arbiter.i_wb_cpu_dbus_dat\[31\] u_scanchain_local.clk u_scanchain_local.module_data_in\[37\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_49_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2302__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2066__B1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__A2 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2823_ _0208_ io_in[4] u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2754_ _0014_ io_in[4] u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1705_ _1136_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2685_ _0074_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1592__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1636_ _1032_ _1024_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1567_ _1014_ _1018_ _1019_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_28_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2541__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1498_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _0960_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1802__C _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2119_ _0467_ _0468_ _0469_ _0470_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1980__S _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2532__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2599__A1 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1646__I0 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[21\]
+ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1421_ _0901_ _0903_ _0906_ u_arbiter.o_wb_cpu_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2806_ _0191_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2737_ _0126_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2668_ _0057_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1619_ _1055_ _1059_ _1062_ u_cpu.cpu.state.stage_two_req _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2599_ u_cpu.cpu.decode.co_ebreak u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\]
+ _1037_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2514__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2514__B2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1975__S _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2806__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2505__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _1189_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[24\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2441__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2522_ u_cpu.cpu.immdec.imm11_7\[2\] _0764_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1547__A2 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2453_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[13\]
+ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2384_ _0694_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1404_ _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3005_ _3005_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2829__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1786__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1943__C1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[47\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[5] u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1465__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1953_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1884_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _1196_ _0252_ _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2505_ _0340_ _0348_ _0398_ _0419_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1940__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2436_ _0726_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2367_ u_arbiter.i_wb_cpu_dbus_adr\[9\] u_arbiter.i_wb_cpu_dbus_adr\[10\] _0678_
+ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2298_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_rdt\[0\] _0899_ _0631_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1456__A1 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2651__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1931__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1998__A2 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[67\] u_scanchain_local.module_data_in\[66\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[29\] u_scanchain_local.clk u_scanchain_local.module_data_in\[67\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_15_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1907__C1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2175__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _0333_ _0541_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2674__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2152_ _0500_ _0496_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2083_ _0354_ _0425_ _0409_ _0437_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1630__C _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[43\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2985_ _2985_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1936_ _0309_ _0310_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1867_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _1196_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_u_scanchain_local.scan_flop\[58\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1798_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _1200_ _1196_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1913__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2419_ _1053_ _0713_ _0714_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1821__B _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1429__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1983__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1601__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2157__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1904__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2099__B _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2697__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2093__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_A[4] u_cpu.rf_ram.addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1691__I1 u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2770_ _0156_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1721_ u_cpu.rf_ram_if.rdata0\[5\] _1135_ u_cpu.rf_ram_if.rtrig0 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1652_ _1102_ u_cpu.cpu.ctrl.i_iscomp _1041_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1583_ u_cpu.cpu.decode.op22 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2204_ _0426_ _0420_ _0367_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1659__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2135_ _0352_ _0375_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2320__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2066_ _0364_ _0422_ _0405_ _0350_ _0423_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2084__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2968_ _2968_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1919_ _0298_ _0299_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2899_ _2899_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2311__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1978__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2075__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1822__A1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1889__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2302__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2712__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2066__B2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1664__I1 u_cpu.rf_ram.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2822_ _0207_ io_in[4] u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2753_ _0142_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ u_cpu.rf_ram_if.rdata1\[4\] _1135_ _1010_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2684_ _0073_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1635_ _1032_ _1024_ u_cpu.cpu.bne_or_bge _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1566_ _1014_ u_cpu.cpu.immdec.imm31 _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1497_ _0907_ _0963_ _0964_ u_arbiter.o_wb_cpu_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2118_ _0367_ _0368_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2049_ _0345_ _0347_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1804__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2735__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2296__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1646__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2599__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2220__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1420_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2523__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2287__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2039__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2805_ _0190_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2736_ _0125_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2667_ _0056_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1565__A3 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1618_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2598_ u_cpu.cpu.genblk3.csr.mie_mtie _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2514__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1549_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2758__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2202__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2505__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2521_ u_cpu.cpu.immdec.imm11_7\[3\] _0382_ _0395_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2452_ _0734_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2383_ u_arbiter.i_wb_cpu_dbus_adr\[17\] u_arbiter.i_wb_cpu_dbus_adr\[18\] _0678_
+ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1403_ io_in[1] _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3004_ _3004_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1483__A2 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2719_ _0108_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1943__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2499__A1 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2423__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1785__I _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1777__A3 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[12\] u_arbiter.i_wb_cpu_rdt\[9\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA_u_cpu.rf_ram.RAM0_D[4] u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2284__C _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1952_ _0320_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1883_ _1196_ _1197_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2504_ _1015_ _0764_ _0765_ _0601_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2435_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[4\]
+ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2366_ _0685_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2297_ _0615_ _0607_ _0629_ _0630_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[10\]_D u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1392__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[14\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1447__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[8\]_D u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1907__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2220_ _0421_ _0561_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2819__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2151_ u_cpu.cpu.immdec.imm24_20\[1\] _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2082_ _0343_ _0388_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_47_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2984_ _2984_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ u_arbiter.i_wb_cpu_rdt\[19\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1866_ _0254_ _0255_ _0259_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1797_ _1014_ _1061_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[37\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2418_ u_cpu.cpu.bufreg.lsb\[1\] _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2349_ _0674_ _0675_ _0676_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1601__A2 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_scanchain_local.scan_flop\[5\] u_arbiter.i_wb_cpu_rdt\[2\] io_in[3] u_arbiter.i_wb_cpu_dbus_sel\[3\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2617__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2093__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_cpu.rf_ram.RAM0_A[3] u_cpu.rf_ram.addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1840__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1720_ _1145_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1651_ u_cpu.cpu.state.o_cnt_r\[2\] u_cpu.cpu.ctrl.i_iscomp _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2070__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2641__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1582_ _1012_ _1013_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2203_ _0354_ _0370_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2134_ _0343_ _0375_ _0371_ _0370_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_6_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2791__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2608__A1 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2065_ _0857_ _1192_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2967_ _2967_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2898_ _2898_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1918_ u_arbiter.i_wb_cpu_rdt\[13\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1595__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1849_ _1016_ _0245_ _0032_ _0857_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1822__A2 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1994__S _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2664__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1586__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1889__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[42\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[57\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2821_ _0206_ io_in[4] u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2752_ _0141_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1703_ _1128_ _0021_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2683_ _0072_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1634_ _0860_ _1032_ _1024_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1565_ _0855_ u_cpu.cpu.branch_op _0853_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1496_ u_arbiter.i_wb_cpu_dbus_adr\[20\] _0926_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1652__B _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1501__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2117_ _0448_ _0458_ _0369_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2057__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2048_ _1192_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2687__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1804__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1568__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2296__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1646__I2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2599__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[42\] u_scanchain_local.module_data_in\[41\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[4\] u_scanchain_local.clk u_scanchain_local.module_data_in\[42\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_6_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2039__A2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2804_ _0189_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2735_ _0124_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2666_ _0055_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1970__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1617_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2597_ _0830_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1548_ _0858_ _0861_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1479_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _0949_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1789__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2702__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2852__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2441__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2520_ _0379_ _0776_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2451_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[12\]
+ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1402_ _0851_ u_cpu.rf_ram_if.wtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_64_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2382_ _0693_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3003_ _3003_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1483__A3 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2725__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2718_ _0107_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1943__A1 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2649_ _0038_ io_in[4] u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1777__A4 u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2187__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[3] u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2111__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2748__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1951_ u_arbiter.i_wb_cpu_rdt\[25\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2414__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1882_ _0257_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2178__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2503_ u_cpu.cpu.immdec.imm11_7\[1\] _0334_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2434_ _0725_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_9_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2365_ u_arbiter.i_wb_cpu_dbus_adr\[8\] u_arbiter.i_wb_cpu_dbus_adr\[9\] _0678_ _0685_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2296_ u_cpu.cpu.immdec.imm19_12_20\[5\] _0334_ _0607_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2102__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1392__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2341__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2158__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1907__A1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2332__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ _0495_ _0498_ _0499_ _0455_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2081_ _0336_ _0350_ _0411_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2983_ _2983_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_59_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1934_ u_arbiter.i_wb_cpu_dbus_dat\[20\] _0286_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1865_ u_arbiter.i_wb_cpu_rdt\[0\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1796_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2417_ _1064_ _1195_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2348_ u_cpu.cpu.genblk3.csr.mie_mtie u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.i_mtip
+ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2279_ u_cpu.cpu.csr_imm _0334_ _0606_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2827__D _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2093__A3 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[2] u_cpu.rf_ram.addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1650_ u_cpu.cpu.state.o_cnt_r\[1\] _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1581_ _1031_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2305__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2202_ _0494_ _0545_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2133_ _0457_ _0481_ _0483_ _0479_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2064_ _0345_ _0420_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2608__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2966_ _2966_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2897_ _2897_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1917_ u_arbiter.i_wb_cpu_dbus_dat\[14\] _0286_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2092__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1595__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1848_ u_cpu.cpu.bne_or_bge _0244_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1779_ u_cpu.cpu.immdec.imm11_7\[4\] _1185_ _1186_ _1181_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[11\]_SI u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1404__I _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2480__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2809__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1586__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2535__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[27\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ _0205_ io_in[4] u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2751_ _0140_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2682_ _0071_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1702_ _1134_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ _0866_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2526__A1 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1564_ u_arbiter.i_wb_cpu_dbus_we _1017_ u_cpu.cpu.immdec.imm24_20\[0\] _1019_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1495_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _0960_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2116_ _0369_ _0448_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2047_ _0396_ _0400_ _0406_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2462__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2949_ _2949_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1568__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2517__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1740__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1646__I3 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2453__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2599__A4 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2781__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[35\] u_scanchain_local.module_data_in\[34\] io_in[3]
+ u_arbiter.i_wb_cpu_dbus_dat\[29\] u_scanchain_local.clk u_scanchain_local.module_data_in\[35\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1495__A1 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2141__C1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1798__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2803_ _0188_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2734_ _0123_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2665_ _0054_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1970__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2596_ u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.mstatus_mpie _0829_
+ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1616_ _1017_ _1067_ _1068_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ u_arbiter.i_wb_cpu_dbus_we u_cpu.cpu.bufreg.i_sh_signed _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1478_ _0905_ _0947_ _0949_ _0950_ u_arbiter.o_wb_cpu_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_41_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2654__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2435__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[41\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[56\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__A4 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2450_ _0733_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1401_ _0880_ _0890_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2381_ u_arbiter.i_wb_cpu_dbus_adr\[16\] u_arbiter.i_wb_cpu_dbus_adr\[17\] _0678_
+ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2677__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3002_ _3002_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1640__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2717_ _0106_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1943__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2648_ _0037_ io_in[4] u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2579_ _1014_ _0873_ _1045_ _1038_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1412__I _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1631__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2187__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1934__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[2] u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2111__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1870__A1 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ _0318_ _0319_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1881_ u_arbiter.i_wb_cpu_rdt\[3\] _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2502_ _1192_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2433_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[3\]
+ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2102__B _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2364_ _0684_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2295_ _0407_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2102__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1861__A1 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1613__A1 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2842__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2169__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2341__A2 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[60\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1907__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2332__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2080_ _0424_ _0407_ _0436_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2096__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2715__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__B _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2982_ _2982_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1933_ _0307_ _0308_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1864_ _0257_ _0252_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1795_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2416_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] _1038_ _1195_ _0712_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2347_ _1014_ _1181_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2278_ u_cpu.cpu.immdec.imm19_12_20\[3\] _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2087__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1834__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2738__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[8\]_SI u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2078__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[1] u_cpu.rf_ram.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1825__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1600__I _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[65\] u_scanchain_local.module_data_in\[64\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[27\] u_scanchain_local.clk u_scanchain_local.module_data_in\[65\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2250__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2002__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1580_ _0853_ _1032_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2201_ u_cpu.cpu.immdec.imm30_25\[1\] _0542_ _0544_ u_cpu.cpu.immdec.imm30_25\[2\]
+ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2132_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2063_ _1192_ _0404_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1816__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2965_ _2965_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2896_ _2896_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1916_ _0297_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2092__I1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1847_ _0238_ _0242_ _0243_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1778_ _1016_ u_arbiter.i_wb_cpu_dbus_we _1107_ _0856_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2232__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1586__A3 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2535__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2299__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2838__D u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2750_ _0139_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2223__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2681_ _0070_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1701_ u_cpu.rf_ram_if.rdata1\[3\] _1133_ _1010_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1632_ _1084_ _1003_ _1024_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1563_ u_arbiter.i_wb_cpu_dbus_we _1015_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1494_ _0905_ _0960_ _0961_ _0962_ u_arbiter.o_wb_cpu_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2110__B _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2115_ _1189_ u_arbiter.i_wb_cpu_rdt\[4\] _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2046_ _0855_ _0334_ _0355_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2462__A1 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2948_ _2948_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2214__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2879_ _2879_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2517__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1740__A3 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1964__B1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2508__A2 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[28\] u_arbiter.i_wb_cpu_rdt\[25\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1495__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2141__C2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2357__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2802_ _0187_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2092__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2733_ _0122_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2664_ _0053_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2595_ _1014_ _0873_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1615_ _1016_ u_cpu.cpu.decode.opcode\[1\] _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1546_ _1001_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_8_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1477_ u_arbiter.i_wb_cpu_dbus_adr\[15\] _0926_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2029_ u_cpu.cpu.decode.opcode\[1\] _0334_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1946__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[17\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1477__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2426__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2851__D u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[31\]_D u_arbiter.i_wb_cpu_rdt\[28\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1400_ _0884_ _0885_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_64_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2380_ _0692_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3001_ _3001_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1468__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2417__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[22\]_D u_arbiter.i_wb_cpu_rdt\[19\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_2716_ _0105_ io_in[4] u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2647_ _0036_ io_in[4] u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2578_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _0816_ _0872_ _0817_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1529_ _0907_ _0987_ _0988_ u_arbiter.o_wb_cpu_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1459__A2 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2771__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[13\]_D u_arbiter.i_wb_cpu_rdt\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2344__B1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_cpu.rf_ram.RAM0_D[1] u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2846__D u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1880_ _0271_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1622__A2 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1386__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2501_ _1165_ _1186_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2432_ _0724_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_116_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2363_ u_arbiter.i_wb_cpu_dbus_adr\[7\] u_arbiter.i_wb_cpu_dbus_adr\[8\] _0678_ _0684_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2794__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2294_ _0397_ _0403_ _0618_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[40\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2545__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[55\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1613__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1392__A4 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2341__A3 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1604__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2667__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2317__B1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[10\] u_arbiter.i_wb_cpu_rdt\[7\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_113_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1540__A1 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2365__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1843__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2981_ _2981_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_43_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1932_ u_arbiter.i_wb_cpu_rdt\[18\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1863_ _0256_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1794_ u_arbiter.i_wb_cpu_dbus_dat\[3\] u_arbiter.i_wb_cpu_dbus_dat\[2\] u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ u_arbiter.i_wb_cpu_dbus_dat\[1\] _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2415_ _0707_ _0709_ _0711_ _1064_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2346_ u_cpu.cpu.genblk3.csr.timer_irq_r _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2277_ _0611_ _0607_ _0612_ _0441_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2087__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1598__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_cpu.rf_ram.RAM0_A[0] u_cpu.rf_ram.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1589__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[58\] u_scanchain_local.module_data_in\[57\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[20\] u_scanchain_local.clk u_scanchain_local.module_data_in\[58\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2002__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1772__B _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2200_ _1192_ _0538_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1513__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2561__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2131_ _0335_ _0413_ _0342_ _0409_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_26_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2062_ _0377_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2832__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2964_ _2964_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1915_ u_arbiter.i_wb_cpu_rdt\[12\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[13\] _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2895_ _2895_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_72_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1846_ u_cpu.cpu.alu.cmp_r _1091_ _1085_ _0238_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1777_ u_cpu.cpu.immdec.imm11_7\[1\] u_cpu.cpu.immdec.imm11_7\[2\] u_cpu.cpu.immdec.imm11_7\[3\]
+ u_cpu.cpu.immdec.imm11_7\[0\] _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1752__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[50\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2329_ u_cpu.cpu.immdec.imm19_12_20\[8\] _1192_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2480__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1586__A4 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1991__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2705__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2855__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[3\] u_arbiter.i_wb_cpu_rdt\[0\] io_in[3] u_arbiter.i_wb_cpu_dbus_sel\[1\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_64_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2854__D u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2223__A2 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2680_ _0069_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1700_ _1128_ _0020_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1631_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1562_ _0855_ _1016_ u_cpu.cpu.decode.opcode\[1\] _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1493_ u_arbiter.i_wb_cpu_dbus_adr\[19\] _0904_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2114_ _0899_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2045_ _0333_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2553__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2462__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2947_ _2947_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2214__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2728__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2352__I _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2878_ _2878_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1829_ _0230_ _1206_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2517__A3 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2301__B _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2141__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2141__B2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2373__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2801_ _0186_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2732_ _0121_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1955__A1 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2663_ _0052_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1717__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2594_ _0826_ _0827_ _0828_ _1051_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1614_ _0857_ u_arbiter.i_wb_cpu_dbus_we _0863_ _0870_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1545_ _0999_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1476_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _0937_ _0948_
+ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_132_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2028_ _0369_ _0388_ _0381_ _0354_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2435__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1946__A1 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2123__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2426__A2 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_scanchain_local.scan_flop\[40\] u_scanchain_local.module_data_in\[39\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[2\] u_scanchain_local.clk u_scanchain_local.module_data_in\[40\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1780__B _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2114__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3000_ _3000_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2417__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2715_ _0104_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2646_ _0035_ io_in[4] u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2577_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1528_ u_arbiter.i_wb_cpu_dbus_adr\[28\] _0926_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1459_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] u_cpu.cpu.ctrl.o_ibus_adr\[10\] _0936_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2105__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1849__C _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1395__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2344__B2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_D[0] u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1775__B _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2500_ _0891_ _1182_ _0761_ _0762_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_31_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2431_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2335__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2362_ _0683_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2293_ _0619_ _0595_ _0626_ _0338_ _0381_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_29_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[1\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2561__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1377__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2326__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2629_ _0031_ io_in[4] u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[14\]_SI u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2317__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2317__B2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1540__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2096__A3 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ _2980_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1931_ u_arbiter.i_wb_cpu_dbus_dat\[19\] _0286_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1862_ u_arbiter.i_wb_cpu_ack _0904_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2381__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2761__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1793_ _1194_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1725__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2414_ _1173_ _1176_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2345_ _0673_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_42_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2276_ u_cpu.cpu.immdec.imm19_12_20\[3\] _0334_ _0606_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1598__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2634__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2784__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2250__A3 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2538__A1 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[54\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2130_ _0343_ _0385_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[69\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2061_ _0385_ _0361_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2474__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2963_ _2963_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1914_ _0295_ _0296_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2894_ _2894_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_33_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2529__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1845_ _1027_ _0241_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1776_ _0874_ _1165_ u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1752__A2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1504__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2657__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2328_ _0381_ _0654_ _0658_ _0382_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2259_ _0367_ _0590_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1440__A1 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2209__B _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2223__A3 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1630_ _0857_ _1065_ _1082_ _0873_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1982__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1783__B _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1561_ u_cpu.cpu.decode.opcode\[0\] _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1734__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1492_ _0958_ _0959_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1498__A1 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2113_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_rdt\[6\] _0899_ _0465_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2298__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2044_ _0401_ _0402_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2447__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _2946_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2877_ _2877_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ u_cpu.rf_ram_if.rgnt _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1759_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.bufreg.c_r _1168_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_11_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__C _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2150__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1868__B _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1964__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2822__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2141__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2429__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2800_ _0185_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[40\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2731_ _0120_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1955__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ _0051_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.output_buffers\[2\] u_scanchain_local.data_out_i u_scanchain_local.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2593_ u_cpu.cpu.genblk3.csr.o_new_irq _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1613_ u_cpu.cpu.state.o_cnt_r\[0\] _1038_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1544_ u_cpu.rf_ram_if.rcnt\[0\] _0849_ _0850_ u_cpu.rf_ram_if.wen0_r _1000_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1475_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] u_cpu.cpu.ctrl.o_ibus_adr\[14\] _0948_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1891__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ _0385_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2929_ _2929_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2845__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1946__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[63\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1634__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1937__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1617__I _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[33\] u_arbiter.i_wb_cpu_rdt\[30\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_64_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2718__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1625__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1928__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2714_ _0103_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2645_ _0034_ io_in[4] u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2559__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2576_ _0815_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1527_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1458_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _0930_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _0935_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2105__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1864__A1 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1389_ u_cpu.cpu.immdec.imm19_12_20\[8\] _0851_ _0876_ u_cpu.cpu.immdec.imm24_20\[4\]
+ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2344__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1855__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__I0 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2032__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2583__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2430_ _0723_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_68_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2379__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2361_ u_arbiter.i_wb_cpu_dbus_adr\[6\] u_arbiter.i_wb_cpu_dbus_adr\[7\] _0678_ _0683_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2292_ _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2099__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2690__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2271__B2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2326__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2628_ _0030_ io_in[4] u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2559_ u_arbiter.i_wb_cpu_rdt\[23\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _0799_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1837__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2262__B2 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2262__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2317__A2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1930_ _0305_ _0306_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2253__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1861_ u_arbiter.i_wb_cpu_dbus_dat\[1\] _1196_ _1204_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2005__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1792_ _1054_ _1058_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2413_ _1173_ _1176_ _1181_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2344_ u_cpu.cpu.immdec.imm31 _0334_ _0405_ _0671_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2275_ u_cpu.cpu.immdec.imm19_12_20\[2\] _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1819__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2304__C _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2281__I u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _1005_ _0407_ _0418_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1360__I _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2962_ _2962_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2226__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1913_ u_arbiter.i_wb_cpu_rdt\[11\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2893_ _2893_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_37_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2529__A2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1844_ _1032_ _1024_ _0240_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1775_ _1183_ _1184_ _1182_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2567__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2327_ _0360_ _0402_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2258_ _0592_ _0593_ _0594_ _0596_ _0408_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2189_ u_arbiter.i_wb_cpu_rdt\[25\] u_arbiter.i_wb_cpu_rdt\[9\] _0900_ _0534_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1440__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1900__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2751__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[63\] u_scanchain_local.module_data_in\[62\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[25\] u_scanchain_local.clk u_scanchain_local.module_data_in\[63\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1967__B1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1431__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1560_ u_cpu.cpu.immdec.imm11_7\[0\] _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1491_ _0958_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1498__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2387__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2112_ _0864_ _0407_ _0464_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2298__I1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2043_ _0367_ _0347_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2447__B2 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2945_ _2945_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2876_ _2876_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ u_cpu.cpu.state.o_cnt_r\[3\] _0228_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1758_ _0857_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1689_ _1125_ u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2774__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[53\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1949__B1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[68\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1884__B _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2429__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2429__B2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__C _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1652__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[34\]_D u_arbiter.i_wb_cpu_rdt\[31\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ _0119_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2661_ _0050_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2647__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1612_ _1053_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2592_ _1014_ _1044_ _0873_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2797__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1543_ u_cpu.rf_ram_if.wen1_r _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1474_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _0942_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _0947_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1891__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2026_ _1189_ u_arbiter.i_wb_cpu_rdt\[13\] _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[25\]_D u_arbiter.i_wb_cpu_rdt\[22\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ _2928_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2580__S _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2859_ _2859_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_123_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[16\]_D u_arbiter.i_wb_cpu_rdt\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1398__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[26\] u_arbiter.i_wb_cpu_rdt\[23\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1789__B _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1625__A2 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1389__B2 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2050__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2413__B _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2713_ _0102_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2189__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2644_ _0033_ io_in[4] u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2575_ u_arbiter.i_wb_cpu_rdt\[31\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _0799_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1526_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] u_cpu.cpu.ctrl.o_ibus_adr\[26\] _0980_ _0986_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1457_ _0932_ _0934_ u_arbiter.o_wb_cpu_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1388_ u_cpu.rf_ram_if.rtrig0 _0875_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2575__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1864__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2113__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2812__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2009_ u_arbiter.i_wb_cpu_rdt\[13\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _0898_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[30\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1855__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2280__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__I1 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2032__A2 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2360_ _0682_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2291_ _0621_ _0622_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2099__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2395__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2835__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1846__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2271__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2627_ _0029_ io_in[4] u_cpu.rf_ram_if.rcnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[53\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2558_ _0806_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1509_ _0907_ _0972_ _0973_ u_arbiter.o_wb_cpu_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2489_ _0753_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_43_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1837__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2014__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2708__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1773__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1525__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2573__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2253__A2 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1860_ _0252_ _0253_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2005__A2 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1791_ _1031_ _0855_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1764__A1 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2412_ u_cpu.cpu.bufreg.i_sh_signed _1181_ _1064_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2343_ _0616_ _0571_ _0480_ _0382_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2274_ _0609_ _0607_ _0610_ _0436_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1755__A1 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2601__B _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2555__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2680__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2171__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2474__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2961_ _2961_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2226__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1912_ u_arbiter.i_wb_cpu_dbus_dat\[12\] _0286_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2892_ _2892_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_72_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1985__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ _1032_ _1024_ _0239_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1737__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1774_ _1104_ _1105_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2162__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2326_ _0336_ _0624_ _0655_ _0656_ _0402_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2257_ _0338_ _0409_ _0595_ _0397_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2188_ _0368_ _0399_ _0532_ _0381_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1728__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1662__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1900__A1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2208__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[56\] u_scanchain_local.module_data_in\[55\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[18\] u_scanchain_local.clk u_scanchain_local.module_data_in\[56\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_32_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1490_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] u_cpu.cpu.ctrl.o_ibus_adr\[17\] u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _0949_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2111_ _0405_ _0456_ _0461_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2042_ _0345_ _0368_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2447__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2416__B _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2944_ _2944_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2875_ _2875_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_31_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _0891_ _1014_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1757_ _1016_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1546__I _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1688_ u_cpu.rf_ram_if.wdata0_r\[6\] u_cpu.rf_ram_if.wdata1_r\[6\] _0998_ _1125_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2135__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2309_ _0632_ _0633_ _0381_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1949__A1 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2126__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[1\] u_cpu.cpu.genblk3.csr.i_mtip io_in[3] u_arbiter.o_wb_cpu_we
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_92_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2429__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2236__B _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2660_ _0049_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1611_ _1060_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2591_ u_cpu.cpu.genblk3.csr.mcause31 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1366__I _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1542_ u_cpu.rf_ram_if.genblk1.wtrig0_r _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1473_ _0944_ _0946_ u_arbiter.o_wb_cpu_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2117__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2025_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_u_scanchain_local.scan_flop\[4\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2146__B _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2927_ _2927_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2858_ _2858_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_102_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2789_ _0175_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2741__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1809_ u_cpu.raddr\[0\] _0216_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2108__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1634__A3 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2595__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2347__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[19\] u_arbiter.i_wb_cpu_rdt\[16\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1570__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1389__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2764__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2712_ _0101_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2643_ _0032_ io_in[4] u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2338__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2189__I1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2574_ _0814_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1525_ _0907_ _0984_ _0985_ u_arbiter.o_wb_cpu_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[52\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1456_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _0930_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1387_ u_cpu.cpu.immdec.imm19_12_20\[7\] _0851_ _0876_ u_cpu.cpu.immdec.imm24_20\[3\]
+ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2510__B2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2361__I1 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[67\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2113__I1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2008_ _0360_ _0361_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1670__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2637__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2501__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2787__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2006__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1791__A2 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1543__A2 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2290_ _0358_ _0623_ _0470_ _0385_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__B _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2626_ _0028_ io_in[4] u_cpu.rf_ram_if.rcnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2557_ u_arbiter.i_wb_cpu_rdt\[22\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _0799_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1508_ u_arbiter.i_wb_cpu_dbus_adr\[23\] _0926_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2488_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[30\]
+ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1439_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _0917_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2334__B _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2486__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _0891_ _1193_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1575__S _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1764__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2802__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _0707_ _1064_ _0708_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1516__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2342_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_rdt\[15\] _0900_ _0671_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2273_ u_cpu.cpu.immdec.imm19_12_20\[2\] _0334_ _0607_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2138__C _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2492__A3 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[20\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1988_ _1189_ u_arbiter.i_wb_cpu_rdt\[6\] _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1755__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2609_ _0421_ _0839_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2468__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2064__B _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2825__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2171__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2960_ _2960_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_43_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2891_ _2891_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1911_ _0293_ _0294_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[43\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1985__A2 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1842_ u_cpu.cpu.bne_or_bge _0853_ _0860_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1737__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1773_ u_arbiter.i_wb_cpu_ibus_adr\[0\] u_cpu.cpu.ctrl.pc_plus_4_cy_r _1183_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2325_ _0413_ _0593_ _0408_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2256_ _0592_ _0385_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2187_ _0343_ _0345_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1425__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2848__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2153__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1900__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[66\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1416__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1967__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[49\] u_scanchain_local.module_data_in\[48\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[11\] u_scanchain_local.clk u_scanchain_local.module_data_in\[49\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2144__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2110_ _0402_ _0462_ _0421_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2041_ _0385_ _0397_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1655__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2943_ _2943_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1407__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2416__C _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2874_ _2874_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_102_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ _0891_ _0227_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1756_ _0857_ u_cpu.cpu.decode.opcode\[1\] _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1687_ _1124_ u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2135__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2308_ _0637_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2239_ _0480_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2670__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2326__C _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1949__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2071__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2126__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1637__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2009__S _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1610_ u_cpu.cpu.state.stage_two_req _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2590_ _0822_ _0818_ _0825_ _1051_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1541_ _0894_ _0996_ _0997_ u_arbiter.o_wb_cpu_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1472_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _0942_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1876__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2693__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2024_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_cpu.rf_ram.RAM0_CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2926_ _2926_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2053__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2857_ u_cpu.cpu.o_wen1 io_in[4] u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1800__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1808_ _1149_ _1207_ _0216_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2788_ _0174_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1739_ _0884_ _0026_ _1157_ _0886_ u_cpu.rf_ram.addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1867__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1668__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2044__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2595__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2347__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.output_buffers\[3\]_I u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2283__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2711_ _0100_ io_in[4] u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2586__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2642_ _0006_ io_in[4] u_cpu.rf_ram_if.rdata0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2573_ u_arbiter.i_wb_cpu_rdt\[30\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _0799_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1524_ u_arbiter.i_wb_cpu_dbus_adr\[27\] _0926_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1455_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _0930_ _0904_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1849__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1386_ _0851_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2007_ _0367_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2274__B2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2026__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2909_ _2909_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_52_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2329__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2501__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2265__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2265__B2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2017__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[31\] u_arbiter.i_wb_cpu_rdt\[28\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2731__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2008__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _0027_ io_in[4] u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2556_ _0805_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1507_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2487_ _0752_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_130_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1438_ _0916_ _0918_ _0919_ u_arbiter.o_wb_cpu_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1369_ _0856_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1470__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2754__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2238__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[51\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1461__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2410__A1 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[66\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2410_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _1064_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2174__B1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2341_ _0607_ _0666_ _0669_ _0670_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1921__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2272_ u_cpu.cpu.immdec.imm19_12_20\[1\] _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2229__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[19\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1452__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1987_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2627__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2608_ u_cpu.cpu.ctrl.i_iscomp _0334_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2777__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2539_ u_cpu.cpu.bufreg.i_sh_signed _0334_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2468__B2 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1676__S _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2080__B _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[4\]_D u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2890_ _2890_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_76_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1910_ u_arbiter.i_wb_cpu_rdt\[10\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1434__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1841_ _0860_ _0853_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1772_ _1178_ _1180_ _1182_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1993__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1737__A3 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2324_ _0370_ _0388_ _0449_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2255_ _0343_ _0393_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2186_ _0345_ _0528_ _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2165__B _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2138__B1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2075__B _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1975__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _0344_ _0347_ _0398_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_78_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[10\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1655__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2942_ _2942_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1407__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2604__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2873_ _2873_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2080__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1824_ u_cpu.cpu.mem_bytecnt\[1\] _0226_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1755_ _1005_ _0894_ u_arbiter.o_wb_cpu_we vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1591__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1686_ u_cpu.rf_ram_if.wdata0_r\[5\] u_cpu.rf_ram_if.wdata1_r\[5\] _0998_ _1124_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2307_ _0379_ _0399_ _0639_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2238_ _0340_ _0388_ _0570_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2815__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2169_ u_cpu.cpu.immdec.imm24_20\[3\] _0498_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[28\]_D u_arbiter.i_wb_cpu_rdt\[25\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2071__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1582__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[33\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[19\]_D u_arbiter.i_wb_cpu_rdt\[16\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2062__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[61\] u_scanchain_local.module_data_in\[60\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[23\] u_scanchain_local.clk u_scanchain_local.module_data_in\[61\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1540_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _0894_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1573__A1 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1471_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _0942_ _0904_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2838__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2373__I0 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2494__I _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2023_ u_arbiter.i_wb_cpu_rdt\[14\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _0898_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2925_ _2925_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2856_ u_cpu.cpu.o_wen0 io_in[4] u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1800__A2 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1807_ _0215_ _0849_ _0850_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2787_ _0173_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[56\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1738_ u_cpu.cpu.immdec.imm11_7\[1\] _1126_ _0026_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1564__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1669_ _1115_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1867__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2044__A2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1684__S _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2035__A2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2263__B _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ _0099_ io_in[4] u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2641_ _0005_ io_in[4] u_cpu.rf_ram_if.rdata0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2660__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2572_ _0813_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1523_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1454_ u_arbiter.i_wb_cpu_dbus_adr\[10\] _0905_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1385_ _0862_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2006_ u_arbiter.i_wb_cpu_rdt\[1\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _0899_
+ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2274__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2026__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2908_ _2908_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_104_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2839_ u_cpu.rf_ram_if.wdata0_r\[5\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1537__A1 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2017__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2683__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[24\] u_arbiter.i_wb_cpu_rdt\[21\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_68_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1700__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2256__A2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2008__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2624_ _1206_ _0848_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2567__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2555_ u_arbiter.i_wb_cpu_rdt\[21\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _0799_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2192__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2486_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[29\]
+ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1506_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] u_cpu.cpu.ctrl.o_ibus_adr\[21\] u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _0960_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_130_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1437_ u_arbiter.i_wb_cpu_dbus_adr\[6\] _0905_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1368_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1758__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2183__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2486__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2238__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1997__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2410__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2260__C _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2174__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2340_ u_cpu.cpu.immdec.imm19_12_20\[8\] _0607_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2174__B2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1921__A1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2271_ _0582_ _0607_ _0608_ _0455_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1988__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ _0345_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2165__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2607_ _0835_ _0836_ _0837_ _0838_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2538_ _1162_ _0764_ _0795_ _0523_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2469_ _0743_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2468__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1979__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2721__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1840_ u_cpu.cpu.ctrl.i_jump _0228_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ _1029_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2147__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2323_ u_arbiter.i_wb_cpu_rdt\[18\] u_arbiter.i_wb_cpu_rdt\[2\] _0900_ _0654_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2254_ _0371_ _0491_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[7\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2185_ _0343_ _0529_ _0482_ _0448_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_55_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2083__B1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2744__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1969_ _0329_ _0282_ _0286_ _1024_ _0331_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2401__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2138__B2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2138__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[50\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2310__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[65\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_u_cpu.rf_ram.RAM0_WEN[7] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2074__B1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2129__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[18\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2301__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2941_ _2941_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2767__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2872_ _2872_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_102_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1823_ u_cpu.cpu.mem_bytecnt\[0\] _0224_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1754_ _1164_ _1167_ _0907_ u_arbiter.o_wb_cpu_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1685_ _1123_ u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2020__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2306_ _0340_ _0348_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2237_ _0411_ _0413_ _0442_ _0576_ _0429_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ u_cpu.cpu.immdec.imm24_20\[4\] _1192_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2099_ _0356_ _0393_ _0379_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1582__A2 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2531__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2086__B _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[54\] u_scanchain_local.module_data_in\[53\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[16\] u_scanchain_local.clk u_scanchain_local.module_data_in\[54\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2070__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1573__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1470_ u_arbiter.i_wb_cpu_dbus_adr\[14\] _0905_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2022_ _1169_ _0334_ _0365_ _0383_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2589__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2924_ _2924_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2855_ u_cpu.cpu.o_wdata1 io_in[4] u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1800__A3 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1806_ u_cpu.rf_ram_if.rcnt\[0\] _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2786_ _0172_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2210__B1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1737_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _0998_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1668_ u_cpu.rf_ram.rdata\[4\] u_cpu.rf_ram.data\[4\] _0026_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1599_ _1051_ _1052_ u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2513__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2504__A1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2504__B2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2355__I1 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1794__A2 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0004_ io_in[4] u_cpu.rf_ram_if.rdata0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2805__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2571_ u_arbiter.i_wb_cpu_rdt\[29\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _0799_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1522_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _0980_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1951__C1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1453_ _0905_ _0928_ _0930_ _0931_ u_arbiter.o_wb_cpu_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1384_ _0868_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1623__B _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2005_ _1189_ u_arbiter.i_wb_cpu_rdt\[0\] _0366_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1482__A1 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2907_ _2907_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA_u_scanchain_local.scan_flop\[23\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2431__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2838_ u_cpu.rf_ram_if.wdata0_r\[4\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2769_ _0155_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1537__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[30\]_SI u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2828__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__S _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1776__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1528__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[17\] u_arbiter.i_wb_cpu_rdt\[14\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2258__C _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1700__A2 _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[46\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1464__A1 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2623_ _1193_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2554_ _0804_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2567__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1505_ _0907_ _0969_ _0970_ u_arbiter.o_wb_cpu_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2485_ _0751_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1436_ _0894_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1367_ u_cpu.cpu.branch_op _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1455__A1 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1915__C1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[69\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2650__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2314__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2174__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1921__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2270_ u_cpu.cpu.immdec.imm19_12_20\[1\] _0334_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1988__A2 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1985_ _1189_ u_arbiter.i_wb_cpu_rdt\[1\] _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2606_ u_cpu.cpu.genblk3.csr.mstatus_mie _0829_ _0836_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2165__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2537_ _0793_ _0794_ _0764_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1912__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2468_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1419_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2399_ u_arbiter.i_wb_cpu_dbus_adr\[25\] u_arbiter.i_wb_cpu_dbus_adr\[26\] _1073_
+ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2673__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1428__A1 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1979__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1443__A4 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1973__S _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2156__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1770_ _1054_ _1058_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2147__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2322_ _0607_ _0651_ _0652_ _0653_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2696__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2253_ _1189_ u_arbiter.i_wb_cpu_rdt\[7\] _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2184_ _0457_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1658__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2083__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1830__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1968_ u_arbiter.i_wb_cpu_rdt\[31\] _1204_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1899_ u_arbiter.i_wb_cpu_dbus_dat\[7\] _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2138__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1649__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_WEN[6] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2074__B2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2074__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1821__A1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1672__I1 u_cpu.rf_ram.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2129__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1888__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2940_ _2940_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2065__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2871_ _2871_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__1677__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1822_ u_cpu.cpu.mem_bytecnt\[0\] _0224_ _0225_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1753_ u_cpu.cpu.state.init_done _1165_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ u_cpu.rf_ram_if.wdata0_r\[4\] u_cpu.rf_ram_if.wdata1_r\[4\] _0998_ _1123_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1879__A1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2305_ _0358_ _0623_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2236_ _0413_ _0343_ _0411_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2167_ _0381_ _0505_ _0513_ _0382_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2098_ _0344_ _0363_ _0451_ _0356_ _0347_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2056__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2711__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1803__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2516__C1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2295__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1698__S _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[47\] u_scanchain_local.module_data_in\[46\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[9\] u_scanchain_local.clk u_scanchain_local.module_data_in\[47\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1573__A3 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_scanchain_local.input_buf_clk_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2021_ _0369_ _0378_ _0381_ _0356_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_36_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2734__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2286__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2589__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2923_ _2923_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2854_ u_cpu.rf_ram_if.wdata1_r\[7\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2785_ _0171_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1805_ u_cpu.rf_ram_if.rcnt\[0\] _1207_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2210__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1736_ _0889_ _1001_ _1154_ _1155_ u_cpu.rf_ram.addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[64\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1667_ _1114_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1598_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _0873_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2219_ _0480_ _0558_ _0560_ _0379_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_45_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2277__B2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2407__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2029__A1 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[17\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2757__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2268__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1794__A3 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2570_ _0812_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1521_ _0907_ _0981_ _0982_ u_arbiter.o_wb_cpu_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1951__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1452_ u_arbiter.i_wb_cpu_dbus_adr\[9\] _0926_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1383_ _0869_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1690__I _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2259__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _0898_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1482__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2906_ _2906_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_52_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2431__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2837_ u_cpu.rf_ram_if.wdata0_r\[3\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2768_ _0154_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1719_ u_cpu.rf_ram_if.rdata0\[4\] _1133_ u_cpu.rf_ram_if.rtrig0 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2699_ _0088_ io_in[4] u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2498__B2 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1976__S _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1464__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2622_ _0845_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2553_ u_arbiter.i_wb_cpu_rdt\[20\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _0799_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1504_ u_arbiter.i_wb_cpu_dbus_adr\[22\] _0926_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1924__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2484_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[28\]
+ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1435_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\] _0913_ _0917_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1366_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_GWEN _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1915__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1915__C2 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1694__A2 _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[7\]_D u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1382__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[13\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1437__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1984_ _0899_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_u_scanchain_local.out_flop_CLKN u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2605_ u_cpu.cpu.genblk3.csr.mstatus_mpie _0862_ _0886_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2536_ _0382_ _0411_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2467_ _0742_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1418_ _0892_ u_cpu.cpu.state.ibus_cyc _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2398_ _0701_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2818__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1428__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[36\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1978__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2321_ u_cpu.cpu.immdec.imm19_12_20\[6\] _0607_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2252_ _0899_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2183_ _0356_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1830__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1967_ _0327_ _0282_ _0286_ _0329_ _0330_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_u_scanchain_local.scan_flop\[59\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1898_ _0280_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1594__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1594__B2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2519_ _0621_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2640__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2790__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_WEN[5] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1821__A2 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1585__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2065__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ _2870_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1821_ u_cpu.cpu.mem_bytecnt\[0\] _0224_ _0892_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2663__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1752_ _0855_ _0857_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1683_ _1122_ u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1879__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2304_ _0374_ _0593_ _0634_ _0636_ _0408_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2235_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_rdt\[14\] _0900_ _0575_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2166_ _0379_ _0509_ _0511_ _0512_ _0381_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_54_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2097_ _0385_ _0397_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2999_ _2999_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_cpu.rf_ram.RAM0 u_cpu.rf_ram.RAM0/A[0] u_cpu.rf_ram.RAM0/A[1] u_cpu.rf_ram.RAM0/A[2]
+ u_cpu.rf_ram.RAM0/A[3] u_cpu.rf_ram.RAM0/A[4] u_cpu.rf_ram.RAM0/A[5] u_cpu.rf_ram.RAM0/A[6]
+ u_cpu.rf_ram.RAM0/A[7] u_cpu.rf_ram.RAM0/CEN u_cpu.rf_ram.RAM0/CLK u_cpu.rf_ram.RAM0/D[0]
+ u_cpu.rf_ram.RAM0/D[1] u_cpu.rf_ram.RAM0/D[2] u_cpu.rf_ram.RAM0/D[3] u_cpu.rf_ram.RAM0/D[4]
+ u_cpu.rf_ram.RAM0/D[5] u_cpu.rf_ram.RAM0/D[6] u_cpu.rf_ram.RAM0/D[7] u_cpu.rf_ram.RAM0/GWEN
+ u_cpu.rf_ram.RAM0/Q[0] u_cpu.rf_ram.RAM0/Q[1] u_cpu.rf_ram.RAM0/Q[2] u_cpu.rf_ram.RAM0/Q[3]
+ u_cpu.rf_ram.RAM0/Q[4] u_cpu.rf_ram.RAM0/Q[5] u_cpu.rf_ram.RAM0/Q[6] u_cpu.rf_ram.RAM0/Q[7]
+ u_cpu.rf_ram.RAM0/WEN[0] u_cpu.rf_ram.RAM0/WEN[1] u_cpu.rf_ram.RAM0/WEN[2] u_cpu.rf_ram.RAM0/WEN[3]
+ u_cpu.rf_ram.RAM0/WEN[4] u_cpu.rf_ram.RAM0/WEN[5] u_cpu.rf_ram.RAM0/WEN[6] u_cpu.rf_ram.RAM0/WEN[7]
+ vdd vss gf180mcu_fd_ip_sram__sram256x8m8wm1
XANTENNA__1567__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2516__C2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__B1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2686__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2020_ _0333_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2286__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2038__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2922_ _2922_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__1797__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2853_ u_cpu.rf_ram_if.wdata1_r\[6\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2784_ _0170_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1804_ _1193_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1549__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1735_ u_cpu.cpu.immdec.imm11_7\[0\] _0998_ _0873_ _1001_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_89_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1666_ u_cpu.rf_ram.rdata\[3\] u_cpu.rf_ram.data\[3\] _0026_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1597_ _0886_ _1050_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ _0337_ _0433_ _0559_ _0401_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2277__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2149_ u_cpu.cpu.immdec.imm24_20\[0\] _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2029__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1794__A4 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2132__I _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1520_ u_arbiter.i_wb_cpu_dbus_adr\[26\] _0926_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1951__A1 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1451_ _0929_ _0922_ _0923_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1382_ u_cpu.cpu.genblk3.csr.o_new_irq _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2701__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1703__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2851__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2003_ _0344_ _0364_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_24_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2905_ _2905_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2431__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2836_ u_cpu.rf_ram_if.wdata0_r\[2\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2767_ _0153_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1718_ _1144_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2698_ _0087_ io_in[4] u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1649_ _0853_ _1100_ _0855_ _1016_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_28_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2724__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2186__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2110__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[63\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2413__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2290__C _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2621_ _0215_ u_cpu.rf_ram_if.rcnt\[1\] _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2177__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2552_ _0803_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1924__A1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1503_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2483_ _0750_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1434_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _0913_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _0916_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_u_scanchain_local.scan_flop\[16\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1365_ u_cpu.cpu.decode.opcode\[2\] _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2101__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2747__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2819_ _0204_ io_in[4] u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2168__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1915__A1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1735__B _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[22\] u_arbiter.i_wb_cpu_rdt\[19\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1382__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2331__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1983_ u_arbiter.i_wb_cpu_rdt\[0\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _0899_
+ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2604_ _0755_ _1040_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2535_ _0404_ _0419_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2466_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1417_ _0894_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2397_ u_arbiter.i_wb_cpu_dbus_adr\[24\] u_arbiter.i_wb_cpu_dbus_adr\[25\] _1073_
+ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__I1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2322__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1684__I0 u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2313__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2077__B1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2320_ u_cpu.cpu.immdec.imm19_12_20\[7\] _1192_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2251_ _0368_ _0588_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2182_ _0394_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2296__B _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1966_ u_arbiter.i_wb_cpu_rdt\[30\] _1204_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1897_ _0284_ _0285_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1594__A2 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[9\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _0473_ _0479_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2543__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2449_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[11\]
+ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_WEN[4] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[10\]_SI u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2470__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1820_ _0891_ _0223_ _0224_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2808__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[3\]
+ u_cpu.cpu.state.o_cnt_r\[2\] _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1682_ u_cpu.rf_ram_if.wdata0_r\[3\] u_cpu.rf_ram_if.wdata1_r\[3\] _0998_ _1122_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2303_ _0616_ _0479_ _0551_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2234_ _0405_ _0567_ _0573_ _0395_ _0574_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2165_ _0427_ _0433_ _0379_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1500__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2096_ _0345_ _0447_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_u_scanchain_local.scan_flop\[26\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1803__A3 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2998_ _2998_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1949_ u_arbiter.i_wb_cpu_rdt\[24\] _0257_ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2516__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__B2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[49\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1494__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2293__C _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2921_ _2921_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_91_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2630__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2443__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2852_ u_cpu.rf_ram_if.wdata1_r\[5\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2783_ _0169_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1803_ u_cpu.cpu.state.init_done _0869_ _1165_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_141_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2780__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1734_ _0865_ _0886_ _1126_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1665_ _1113_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1596_ u_cpu.cpu.bne_or_bge _1035_ _1048_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2217_ u_arbiter.i_wb_cpu_rdt\[28\] u_arbiter.i_wb_cpu_rdt\[12\] _0900_ _0559_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1485__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2148_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2079_ _0407_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2653__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1738__B _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[52\] u_scanchain_local.module_data_in\[51\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[14\] u_scanchain_local.clk u_scanchain_local.module_data_in\[52\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1951__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1450_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1381_ u_cpu.cpu.decode.op21 _0870_ _0866_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2002_ _0348_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2904_ _2904_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_32_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ u_cpu.rf_ram_if.wdata0_r\[1\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2195__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2766_ _0152_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1717_ u_cpu.rf_ram_if.rdata0\[3\] _1131_ u_cpu.rf_ram_if.rtrig0 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2697_ _0086_ io_in[4] u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1648_ _1097_ _1098_ _1100_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1579_ _0853_ u_cpu.cpu.csr_imm _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2676__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1458__A1 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1402__I _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1630__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1621__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2620_ u_cpu.rf_ram_if.rcnt\[0\] _0850_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2551_ u_arbiter.i_wb_cpu_rdt\[19\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _0799_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2177__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2482_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1924__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1502_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] u_cpu.cpu.ctrl.o_ibus_adr\[20\] _0960_ _0968_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2699__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1433_ _0907_ _0914_ _0915_ u_arbiter.o_wb_cpu_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1364_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2101__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2818_ _0203_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2749_ _0138_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1892__I _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2168__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1915__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2340__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1851__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1603__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2841__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[15\] u_arbiter.i_wb_cpu_rdt\[12\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_46_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2331__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.input_buf_clk io_in[0] u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_19_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1842__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1982_ _0341_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2603_ _0755_ _1050_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2534_ _0398_ _0379_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2465_ _0741_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2396_ _0700_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1416_ _0900_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2322__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2714__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2048__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2086__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1684__I1 u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2010__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[62\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2313__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2077__B2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2077__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1824__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[15\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _0338_ _0398_ _0419_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2069__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[7\]_SI u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2181_ _0371_ _0375_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2737__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1701__S _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1815__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__I1 u_cpu.rf_ram.data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1965_ u_arbiter.i_wb_cpu_dbus_dat\[31\] _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2240__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1896_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _0258_ _0280_ _1202_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2240__B2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2517_ _0337_ _0394_ _0491_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2448_ _0732_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_116_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2379_ u_arbiter.i_wb_cpu_dbus_adr\[15\] u_arbiter.i_wb_cpu_dbus_adr\[16\] _0678_
+ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2059__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_WEN[3] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2534__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2828__D _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[8\] u_arbiter.i_wb_cpu_rdt\[5\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_48_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2470__A1 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1750_ _1031_ _1163_ _0861_ _1053_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_8_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _1121_ u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2302_ _0340_ _0409_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2233_ u_cpu.cpu.immdec.imm30_25\[4\] _0539_ _0563_ u_cpu.cpu.immdec.imm30_25\[5\]
+ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2289__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2164_ _0385_ _0505_ _0510_ _0491_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2095_ _0438_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1803__A4 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2997_ _2997_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1948_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _0282_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1879_ u_arbiter.i_wb_cpu_rdt\[2\] _1204_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2516__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2204__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1494__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2920_ _2920_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[8\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2851_ u_cpu.rf_ram_if.wdata1_r\[4\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2782_ _0168_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1802_ _0856_ _1203_ _1204_ _0858_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1733_ _1153_ u_cpu.rf_ram.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1664_ u_cpu.rf_ram.rdata\[2\] u_cpu.rf_ram.data\[2\] _0026_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1595_ _0860_ u_cpu.cpu.bne_or_bge _1034_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2216_ _0337_ _0388_ _0393_ _0343_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2147_ _0333_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2078_ _0408_ _0431_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2122__B1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2841__D u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[30\]_D u_arbiter.i_wb_cpu_rdt\[27\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[45\] u_scanchain_local.module_data_in\[44\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[7\] u_scanchain_local.clk u_scanchain_local.module_data_in\[45\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1754__B _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1380_ _0855_ _0857_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[16\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2001_ _0358_ _0362_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2416__A1 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2903_ _2903_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_56_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2834_ _0210_ io_in[4] u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[21\]_D u_arbiter.i_wb_cpu_rdt\[18\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_2765_ _0151_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1716_ _1143_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2696_ _0085_ io_in[4] u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1647_ _1098_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1578_ u_cpu.cpu.alu.i_rs1 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1630__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[12\]_D u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1918__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[39\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1394__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1697__A2 _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2836__D u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2770__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1621__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2550_ _0802_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1385__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2481_ _0749_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1501_ _0907_ _0966_ _0967_ u_arbiter.o_wb_cpu_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1432_ u_arbiter.i_wb_cpu_dbus_adr\[5\] _0905_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1704__S _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1363_ u_cpu.cpu.csr_d_sel _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1999__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1612__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2817_ _0202_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2748_ _0137_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1376__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2643__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2679_ _0068_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2793__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1413__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1851__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1603__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2095__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2582__C _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1842__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2355__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1981_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2666__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2602_ _0831_ _0833_ _0834_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2533_ _0345_ _0451_ _0457_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2158__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2464_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[18\]
+ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2395_ u_arbiter.i_wb_cpu_dbus_adr\[23\] u_arbiter.i_wb_cpu_dbus_adr\[24\] _1073_
+ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1415_ _0900_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3016_ u_scanchain_local.data_out io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2086__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1597__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2010__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1521__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2689__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1588__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1760__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2180_ _0522_ _0525_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2068__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1815__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1964_ _0326_ _0282_ _0286_ _0327_ _0328_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1579__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2240__A2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1895_ u_arbiter.i_wb_cpu_rdt\[5\] _0273_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2516_ _0397_ _0355_ _0393_ _0426_ _0401_ _0337_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_130_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1751__A1 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2447_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[10\]
+ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2551__I0 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2378_ _0691_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1898__I _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2831__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_WEN[2] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1990__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1742__B2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2470__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1680_ u_cpu.rf_ram_if.wdata0_r\[2\] u_cpu.rf_ram_if.wdata1_r\[2\] _0998_ _1121_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2704__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2301_ _0426_ _0375_ _0371_ _0370_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2232_ _0510_ _0568_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2289__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2854__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2163_ _0413_ _0397_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2094_ _0343_ _0425_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[61\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ _2996_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1947_ _0316_ _0317_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1878_ _0266_ _0268_ _1204_ _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[14\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[29\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2727__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1963__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2140__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2443__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2850_ u_cpu.rf_ram_if.wdata1_r\[3\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2363__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1801_ u_arbiter.i_wb_cpu_ack _0904_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2781_ _0167_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1732_ u_cpu.raddr\[1\] _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1663_ _1112_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1707__S _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1706__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1594_ _0868_ _1036_ _1040_ u_cpu.cpu.genblk3.csr.mstatus_mie _1047_ _1048_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2215_ _0484_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_38_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2131__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2146_ _1016_ _1005_ _0859_ _1029_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2077_ _0343_ _0432_ _0433_ _0348_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2979_ _2979_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2198__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1945__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2122__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2122__B2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1476__A3 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[38\] u_scanchain_local.module_data_in\[37\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[0\] u_scanchain_local.clk u_scanchain_local.module_data_in\[38\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_45_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2000_ _0360_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1467__A3 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2902_ _2902_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2416__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2106__B _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2833_ _0025_ io_in[4] u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2764_ _0150_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1715_ u_cpu.rf_ram_if.rdata0\[2\] _1129_ u_cpu.rf_ram_if.rtrig0 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2695_ _0084_ io_in[4] u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1646_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[8\] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_arbiter.i_wb_cpu_dbus_dat\[24\] _0852_ u_cpu.cpu.bufreg.lsb\[1\] _1099_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1577_ _0860_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_28_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2104__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2129_ _0343_ _0479_ _0369_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2067__I u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1918__A1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1918__B2 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1855__B u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1394__A2 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[7\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2343__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2852__D u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2582__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2480_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1500_ u_arbiter.i_wb_cpu_dbus_adr\[21\] _0926_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1431_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2334__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1362_ _0852_ u_cpu.cpu.bufreg.lsb\[1\] u_arbiter.i_wb_cpu_dbus_sel\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2551__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2816_ _0201_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2747_ _0136_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2678_ _0067_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1376__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1629_ _0857_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2325__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[0\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ u_arbiter.i_wb_cpu_rdt\[12\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _0898_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2371__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2601_ _1050_ _0833_ _0892_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2532_ _0407_ _0786_ _0790_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2158__I1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2463_ _0740_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2307__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1715__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2394_ _0699_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1414_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3015_ u_scanchain_local.clk_out io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[29\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2760__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2482__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2204__B _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[20\] u_arbiter.i_wb_cpu_rdt\[17\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1512__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2633__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ u_arbiter.i_wb_cpu_rdt\[29\] _1204_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2783__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1894_ _0281_ _0283_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1579__A2 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2528__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2515_ _0772_ _0775_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1751__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2446_ _0731_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_64_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2377_ u_arbiter.i_wb_cpu_dbus_adr\[14\] u_arbiter.i_wb_cpu_dbus_adr\[15\] _0678_
+ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2464__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_WEN[1] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2216__B1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1990__A2 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1419__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1742__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2656__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2455__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2207__B1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[68\] u_scanchain_local.module_data_in\[67\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[30\] u_scanchain_local.clk u_scanchain_local.module_data_in\[68\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1430__A1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ _0340_ _0385_ _0379_ _0433_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2231_ _0569_ _0571_ _0480_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1497__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2162_ _0427_ _0506_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2093_ _0356_ _0387_ _0419_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2995_ _2995_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1957__C1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1946_ u_arbiter.i_wb_cpu_rdt\[23\] _0273_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _0262_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2679__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2429_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _0719_ _0722_ u_arbiter.i_wb_cpu_ibus_adr\[1\]
+ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2437__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1963__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1479__A1 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2140__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _0860_ _0854_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2780_ _0166_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ u_cpu.raddr\[0\] _1150_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1662_ u_cpu.rf_ram.rdata\[1\] u_cpu.rf_ram.data\[1\] _0026_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2821__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1593_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1723__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2214_ _0467_ _0375_ _0485_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2131__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2145_ u_cpu.cpu.immdec.imm24_20\[1\] _0382_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2076_ _0385_ _0361_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2978_ _2978_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1929_ u_arbiter.i_wb_cpu_rdt\[17\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1945__A2 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2021__C _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2122__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1633__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2844__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[60\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1872__A1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2901_ _2901_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__1624__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[62\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2106__C _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2832_ _0024_ io_in[4] u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2763_ _0149_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[13\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1714_ _1142_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2694_ _0083_ io_in[4] u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1645_ _1031_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\] _0861_ _1098_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_u_scanchain_local.scan_flop\[28\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1576_ _1030_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2549__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2104__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2717__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2128_ _0387_ _0433_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2059_ _0408_ _0416_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1615__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1918__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1855__C _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1871__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1854__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1606__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1909__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2031__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[50\] u_scanchain_local.module_data_in\[49\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[12\] u_scanchain_local.clk u_scanchain_local.module_data_in\[50\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2582__A2 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1430_ _0897_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] u_cpu.cpu.ctrl.o_ibus_adr\[3\] u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_123_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2334__A2 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1361_ u_cpu.cpu.bufreg.lsb\[0\] _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2369__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2098__B2 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2117__B _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2815_ _0200_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2746_ _0135_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2677_ _0066_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1628_ _1066_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1559_ u_cpu.cpu.bufreg2.i_cnt_done _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2089__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2089__B2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2013__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2189__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1827__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2252__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2004__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ _1039_ _0224_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2531_ _0407_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2462_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _0738_ _0721_ u_cpu.cpu.ctrl.o_ibus_adr\[17\]
+ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2307__A2 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2393_ u_arbiter.i_wb_cpu_dbus_adr\[22\] u_arbiter.i_wb_cpu_dbus_adr\[23\] _1073_
+ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1413_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3014_ io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2243__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[6\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2729_ _0118_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2234__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2234__B2 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[13\] u_arbiter.i_wb_cpu_rdt\[10\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ u_arbiter.i_wb_cpu_dbus_dat\[30\] _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2225__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1893_ u_arbiter.i_wb_cpu_rdt\[4\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_18_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2528__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2514_ _0340_ _0405_ _0774_ _0334_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1751__A3 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2445_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2557__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2376_ _0690_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_WEN[0] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2216__B2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2216__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2040__B _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[0\]_D io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2207__B2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2207__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[19\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2230_ _0482_ _0570_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2161_ _0415_ _0507_ _0469_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2377__S _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2092_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_rdt\[4\] _0900_ _0446_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2750__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2994_ _2994_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1945_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _0280_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2125__B _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1957__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ _0252_ _0267_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1980__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2428_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2359_ u_arbiter.i_wb_cpu_dbus_adr\[5\] u_arbiter.i_wb_cpu_dbus_adr\[6\] _0678_ _0682_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[6\] u_arbiter.i_wb_cpu_rdt\[3\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1479__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2773__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1651__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[33\]_D u_arbiter.i_wb_cpu_rdt\[30\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1730_ _1151_ u_cpu.rf_ram.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2600__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1784__B _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1661_ _1006_ _1009_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1592_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _1041_ _1043_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2213_ _0554_ _0555_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2144_ _0477_ _0494_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2075_ _0408_ _0377_ _0404_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[24\]_D u_arbiter.i_wb_cpu_rdt\[21\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2977_ _2977_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1928_ u_arbiter.i_wb_cpu_dbus_dat\[18\] _0286_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1859_ u_arbiter.i_wb_cpu_dbus_dat\[0\] _1196_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2796__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[15\]_D u_arbiter.i_wb_cpu_rdt\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1872__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1779__B _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2900_ _2900_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_56_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2669__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1624__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2831_ _0023_ io_in[4] u_cpu.rf_ram.rdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2762_ _0148_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1388__A1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1713_ u_cpu.rf_ram_if.rdata0\[1\] _1141_ u_cpu.rf_ram_if.rtrig0 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2693_ _0082_ io_in[4] u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2122__C _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1644_ u_cpu.cpu.mem_if.signbit _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1575_ _1003_ _1027_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2565__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2127_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_rdt\[10\] _0899_ _0478_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2058_ _0367_ _0397_ _0352_ _0381_ _0382_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1615__A2 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2040__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1551__A1 u_cpu.rf_ram.data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2811__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2103__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[43\] u_scanchain_local.module_data_in\[42\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[5\] u_scanchain_local.clk u_scanchain_local.module_data_in\[43\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1790__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1360_ _0851_ u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_62_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2342__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2098__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2385__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2184__I _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2270__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2814_ _0199_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _0134_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2022__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2676_ _0065_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1781__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1627_ _1071_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1533__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1558_ u_cpu.rf_ram_if.rdata1\[0\] _1011_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1489_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2834__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[52\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1827__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[27\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2707__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2530_ _0361_ _0379_ _0429_ _0408_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_6_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2461_ _0739_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1412_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2392_ _0698_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2563__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2857__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3013_ io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2243__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ _0117_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1754__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2659_ _0048_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2310__C _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2482__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2545__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2170__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1961_ u_arbiter.i_wb_cpu_dbus_dat\[29\] _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2225__A2 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ _0258_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1984__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ _1159_ _0763_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2444_ _0730_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2375_ u_arbiter.i_wb_cpu_dbus_adr\[13\] u_arbiter.i_wb_cpu_dbus_adr\[14\] _0678_
+ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2464__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2573__S _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2216__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2455__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2207__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1966__A1 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[5\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2143__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2160_ _0343_ _0425_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2091_ _0854_ _0407_ _0445_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2393__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2993_ _2993_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1944_ _0315_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1957__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1875_ u_arbiter.i_wb_cpu_dbus_dat\[2\] u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ _1196_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_31_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1709__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2427_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2134__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2358_ _0681_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1893__B1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2289_ _0343_ _0397_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2437__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1645__B1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1948__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1446__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2125__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_cpu.rf_ram.RAM0_CEN _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2600__A2 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ _1083_ _1111_ u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1591_ _1029_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_4_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2116__A1 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2212_ u_cpu.cpu.immdec.imm30_25\[2\] _0542_ _0544_ u_cpu.cpu.immdec.imm30_25\[3\]
+ _0549_ _0405_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2131__A4 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2143_ _0405_ _0478_ _0490_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2074_ _0356_ _0425_ _0393_ _0371_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2976_ _2976_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ _0304_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_33_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1858_ _1194_ _0251_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1789_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r u_cpu.cpu.state.stage_two_req
+ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2298__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2107__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[3\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1885__B _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1397__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2740__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__C _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2830_ _0022_ io_in[4] u_cpu.rf_ram.rdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2761_ _0147_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1712_ _1006_ _1009_ u_cpu.rf_ram.regzero _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2692_ _0081_ io_in[4] u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1643_ _1078_ _1066_ _1080_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2337__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1574_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2126_ u_cpu.cpu.decode.op26 _0334_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2057_ _0376_ _0394_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2959_ _2959_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2763__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2328__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2500__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2103__I1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2319__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[36\] u_scanchain_local.module_data_in\[35\] io_in[3]
+ u_arbiter.i_wb_cpu_dbus_dat\[30\] u_scanchain_local.clk u_scanchain_local.module_data_in\[36\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1790__A2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2342__I1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2636__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2786__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2813_ _0198_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _0133_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2133__C _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2675_ _0064_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1781__A2 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1626_ _1074_ _1076_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1557_ _1006_ _1009_ u_cpu.rf_ram.regzero _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1488_ _0957_ u_arbiter.o_wb_cpu_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1480__S _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ _0354_ _0393_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2324__B _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1524__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2659__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2460_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _0738_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1411_ u_cpu.cpu.genblk1.align.ctrl_misal _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2391_ u_arbiter.i_wb_cpu_dbus_adr\[21\] u_arbiter.i_wb_cpu_dbus_adr\[22\] _1073_
+ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1364__I _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3012_ io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2476__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2727_ _0116_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2801__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2658_ _0047_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2589_ _0863_ _0871_ _0818_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1609_ _0853_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _1061_ u_cpu.cpu.state.init_done _1062_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1745__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1902__C1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2170__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1960_ _0325_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_42_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1891_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _1196_ _1198_ _0278_ _0280_ _0281_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1433__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2824__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2512_ u_cpu.cpu.immdec.imm11_7\[1\] _0763_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1736__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2443_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2374_ _0689_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2449__B1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[42\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[11\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[26\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2152__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1415__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2847__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1966__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2143__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2090_ _0407_ _0444_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[65\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1798__B _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1654__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2992_ _2992_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1943_ u_arbiter.i_wb_cpu_rdt\[22\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[23\] _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1957__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2206__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1874_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _1196_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2426_ _0891_ _1182_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2134__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2357_ u_arbiter.i_wb_cpu_dbus_adr\[4\] u_arbiter.i_wb_cpu_dbus_adr\[5\] _0678_ _0681_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1893__B2 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1893__A1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2288_ _0397_ _0388_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1645__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1645__B2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__C _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1948__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2332__B _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2125__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1884__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[66\] u_scanchain_local.module_data_in\[65\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[28\] u_scanchain_local.clk u_scanchain_local.module_data_in\[66\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2061__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1590_ _0864_ u_cpu.cpu.decode.co_ebreak _0867_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_4_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2116__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2211_ _0548_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1875__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2142_ _0402_ _0492_ _0421_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2073_ _0414_ _0428_ _0429_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2417__B _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2975_ _2975_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2052__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1926_ u_arbiter.i_wb_cpu_rdt\[16\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[17\] _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_129_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1857_ _1029_ _0249_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1788_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2107__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2409_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2692__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[4\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2043__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1609__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2282__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2760_ _0146_ io_in[4] u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2034__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1711_ _1140_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2691_ _0080_ io_in[4] u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1642_ _1086_ _1090_ _1093_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2399__S _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2337__A2 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1573_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[3\]
+ u_cpu.cpu.state.o_cnt_r\[2\] _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_28_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1848__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2125_ _1037_ _0407_ _0476_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2056_ _0409_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2958_ _2958_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2025__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1909_ u_arbiter.i_wb_cpu_dbus_dat\[11\] _0286_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2889_ _2889_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_68_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2328__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2500__A2 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2319__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[29\] u_arbiter.i_wb_cpu_rdt\[26\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_62_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1650__I u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2255__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2812_ _0197_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2007__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2743_ _0132_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2674_ _0063_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1625_ _0857_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1556_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1487_ u_arbiter.i_wb_cpu_dbus_adr\[18\] _0956_ _0894_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1560__I u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2108_ _0368_ _0459_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2039_ _0367_ _0385_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2730__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2605__B _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2237__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1410_ _0896_ u_arbiter.o_wb_cpu_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2390_ _0697_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3011_ io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2753__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2228__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2726_ _0115_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2657_ _0046_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1608_ _0860_ _0856_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1506__A3 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2588_ _0821_ _0818_ _0824_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1539_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _0993_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2319__C _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2219__B2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1666__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2626__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[3\]_D u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2776__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1902__B1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1902__C2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1969__B1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1890_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2511_ _0407_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2442_ _0729_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2373_ u_arbiter.i_wb_cpu_dbus_adr\[12\] u_arbiter.i_wb_cpu_dbus_adr\[13\] _0678_
+ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2449__A1 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1424__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2649__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2709_ _0098_ io_in[4] u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2799__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1983__I0 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2137__B1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2612__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1974__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[11\] u_arbiter.i_wb_cpu_rdt\[8\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[5\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2991_ _2991_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1942_ _0313_ _0314_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2603__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1873_ _0265_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_122_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2206__I1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2425_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2356_ _0680_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1893__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2287_ _0408_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1645__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[27\]_D u_arbiter.i_wb_cpu_rdt\[24\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1581__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2530__B1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1884__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2814__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2507__C _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1636__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[18\]_D u_arbiter.i_wb_cpu_rdt\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2061__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2523__B _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xu_scanchain_local.scan_flop\[59\] u_scanchain_local.module_data_in\[58\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[21\] u_scanchain_local.clk u_scanchain_local.module_data_in\[59\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2210_ _0402_ _0550_ _0551_ _0552_ _0421_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[32\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2521__B1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1875__A2 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2141_ _0360_ _0427_ _0362_ _0478_ _0491_ _0338_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_2072_ _0401_ _0387_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[10\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2974_ _2974_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[25\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1925_ _0302_ _0303_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2052__A2 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1856_ u_cpu.cpu.bufreg.lsb\[1\] u_cpu.cpu.mem_bytecnt\[1\] _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1787_ _1189_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1563__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2408_ _0706_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2837__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2363__I0 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2339_ _0857_ _0584_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2043__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1674__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[55\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[4\] u_arbiter.i_wb_cpu_rdt\[1\] io_in[3] u_arbiter.i_wb_cpu_dbus_sel\[2\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_49_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2237__C _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1609__A2 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2282__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2034__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2690_ _0079_ io_in[4] u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1710_ u_cpu.rf_ram_if.rdata1\[6\] _1139_ _1010_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1641_ _0856_ _1057_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1572_ _1004_ _1025_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2124_ _0405_ _0465_ _0475_ _0395_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2055_ _0411_ _0413_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2273__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2957_ _2957_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2888_ _2888_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1908_ _0292_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1784__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1839_ _0235_ _0236_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1536__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2500__A3 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2264__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__B _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2575__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2255__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ _0196_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2007__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2742_ _0131_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2682__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2673_ _0062_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1624_ _0855_ _1016_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1555_ u_cpu.rf_ram_if.rtrig1 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2191__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1486_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _0954_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_u_scanchain_local.scan_flop\[3\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2107_ _0367_ _0354_ _0451_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2038_ _0397_ _0358_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_36_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1509__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2113__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2557__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2182__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2237__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1996__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[41\] u_scanchain_local.module_data_in\[40\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[3\] u_scanchain_local.clk u_scanchain_local.module_data_in\[41\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2023__S _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3010_ io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2476__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2228__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1987__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1739__B2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _0114_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2656_ _0045_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1607_ _1055_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2164__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2587_ u_cpu.cpu.genblk3.csr.o_new_irq _0858_ _0818_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__1506__A4 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1538_ _0992_ _0994_ _0995_ u_arbiter.o_wb_cpu_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1469_ _0905_ _0941_ _0942_ _0943_ u_arbiter.o_wb_cpu_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_80_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1682__S _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1902__A1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1969__B2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2510_ _0766_ _0769_ _0770_ _0402_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2441_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _0719_ _0722_ u_cpu.cpu.ctrl.o_ibus_adr\[7\]
+ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2146__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2720__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2372_ _0688_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1605__B _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2449__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1680__I0 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2171__B _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2708_ _0097_ io_in[4] u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2137__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2137__B2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2639_ _0003_ io_in[4] u_cpu.rf_ram_if.rdata0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1896__B1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[6\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2612__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2081__B _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2743__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[19\]_SI u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2128__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2300__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2990_ _2990_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1941_ u_arbiter.i_wb_cpu_rdt\[21\] _0273_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2603__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1872_ u_arbiter.i_wb_cpu_rdt\[1\] _1204_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2119__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ _1029_ _1181_ _0891_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1590__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2355_ u_arbiter.i_wb_cpu_dbus_adr\[3\] u_arbiter.i_wb_cpu_dbus_adr\[4\] _0678_ _0680_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2286_ _0337_ _0479_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2766__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__B2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2046__B1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2521__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1875__A3 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0360_ _0397_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2639__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2071_ _0426_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2789__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2973_ _2973_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1924_ u_arbiter.i_wb_cpu_rdt\[15\] _0273_ _0282_ u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2206__S _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1855_ u_cpu.cpu.bufreg.lsb\[1\] u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\]
+ _0852_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1786_ u_arbiter.i_wb_cpu_ack _0894_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1563__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2407_ u_arbiter.i_wb_cpu_dbus_adr\[29\] u_arbiter.i_wb_cpu_dbus_adr\[30\] _1073_
+ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2512__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2338_ _0382_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2269_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2028__B1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2579__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2579__B2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1626__I0 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2343__C _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2503__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1793__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1640_ _1074_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1571_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2123_ _0379_ _0472_ _0473_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2054_ _1189_ u_arbiter.i_wb_cpu_rdt\[10\] _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2956_ _2956_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2887_ _2887_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1907_ u_arbiter.i_wb_cpu_rdt\[9\] _0257_ _0258_ u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _0280_ u_arbiter.i_wb_cpu_dbus_dat\[10\] _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_11_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1838_ _1164_ _1166_ _0032_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2804__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1769_ _1078_ _1065_ _1179_ _1071_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1749__I u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[22\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2488__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[24\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2529__B _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[39\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2810_ _0195_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2741_ _0130_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2827__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2672_ _0061_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.output_buffers\[3\] u_scanchain_local.clk u_scanchain_local.clk_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_1623_ u_cpu.cpu.mem_bytecnt\[1\] _1075_ _1022_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1554_ _1007_ _1008_ u_cpu.rf_ram.rdata\[0\] _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1485_ _0905_ _0953_ _0954_ _0955_ u_arbiter.o_wb_cpu_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2191__A2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

