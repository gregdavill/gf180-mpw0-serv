// This is the unpowered netlist.
module serv_2 (io_in,
    io_oeb,
    io_out);
 input [4:0] io_in;
 output [4:0] io_oeb;
 output [4:0] io_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire \u_arbiter.i_wb_cpu_ack ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_we ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[0] ;
 wire \u_arbiter.i_wb_cpu_rdt[10] ;
 wire \u_arbiter.i_wb_cpu_rdt[11] ;
 wire \u_arbiter.i_wb_cpu_rdt[12] ;
 wire \u_arbiter.i_wb_cpu_rdt[13] ;
 wire \u_arbiter.i_wb_cpu_rdt[14] ;
 wire \u_arbiter.i_wb_cpu_rdt[15] ;
 wire \u_arbiter.i_wb_cpu_rdt[16] ;
 wire \u_arbiter.i_wb_cpu_rdt[17] ;
 wire \u_arbiter.i_wb_cpu_rdt[18] ;
 wire \u_arbiter.i_wb_cpu_rdt[19] ;
 wire \u_arbiter.i_wb_cpu_rdt[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[20] ;
 wire \u_arbiter.i_wb_cpu_rdt[21] ;
 wire \u_arbiter.i_wb_cpu_rdt[22] ;
 wire \u_arbiter.i_wb_cpu_rdt[23] ;
 wire \u_arbiter.i_wb_cpu_rdt[24] ;
 wire \u_arbiter.i_wb_cpu_rdt[25] ;
 wire \u_arbiter.i_wb_cpu_rdt[26] ;
 wire \u_arbiter.i_wb_cpu_rdt[27] ;
 wire \u_arbiter.i_wb_cpu_rdt[28] ;
 wire \u_arbiter.i_wb_cpu_rdt[29] ;
 wire \u_arbiter.i_wb_cpu_rdt[2] ;
 wire \u_arbiter.i_wb_cpu_rdt[30] ;
 wire \u_arbiter.i_wb_cpu_rdt[31] ;
 wire \u_arbiter.i_wb_cpu_rdt[3] ;
 wire \u_arbiter.i_wb_cpu_rdt[4] ;
 wire \u_arbiter.i_wb_cpu_rdt[5] ;
 wire \u_arbiter.i_wb_cpu_rdt[6] ;
 wire \u_arbiter.i_wb_cpu_rdt[7] ;
 wire \u_arbiter.i_wb_cpu_rdt[8] ;
 wire \u_arbiter.i_wb_cpu_rdt[9] ;
 wire \u_cpu.cpu.alu.add_cy_r ;
 wire \u_cpu.cpu.alu.cmp_r ;
 wire \u_cpu.cpu.alu.i_rs1 ;
 wire \u_cpu.cpu.bne_or_bge ;
 wire \u_cpu.cpu.branch_op ;
 wire \u_cpu.cpu.bufreg.c_r ;
 wire \u_cpu.cpu.bufreg.i_sh_signed ;
 wire \u_cpu.cpu.bufreg.lsb[0] ;
 wire \u_cpu.cpu.bufreg.lsb[1] ;
 wire \u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \u_cpu.cpu.csr_d_sel ;
 wire \u_cpu.cpu.csr_imm ;
 wire \u_cpu.cpu.ctrl.i_iscomp ;
 wire \u_cpu.cpu.ctrl.i_jump ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \u_cpu.cpu.decode.co_ebreak ;
 wire \u_cpu.cpu.decode.co_mem_word ;
 wire \u_cpu.cpu.decode.op21 ;
 wire \u_cpu.cpu.decode.op22 ;
 wire \u_cpu.cpu.decode.op26 ;
 wire \u_cpu.cpu.decode.opcode[0] ;
 wire \u_cpu.cpu.decode.opcode[1] ;
 wire \u_cpu.cpu.decode.opcode[2] ;
 wire \u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \u_cpu.cpu.genblk3.csr.i_mtip ;
 wire \u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \u_cpu.cpu.immdec.imm11_7[0] ;
 wire \u_cpu.cpu.immdec.imm11_7[1] ;
 wire \u_cpu.cpu.immdec.imm11_7[2] ;
 wire \u_cpu.cpu.immdec.imm11_7[3] ;
 wire \u_cpu.cpu.immdec.imm11_7[4] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \u_cpu.cpu.immdec.imm24_20[0] ;
 wire \u_cpu.cpu.immdec.imm24_20[1] ;
 wire \u_cpu.cpu.immdec.imm24_20[2] ;
 wire \u_cpu.cpu.immdec.imm24_20[3] ;
 wire \u_cpu.cpu.immdec.imm24_20[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[0] ;
 wire \u_cpu.cpu.immdec.imm30_25[1] ;
 wire \u_cpu.cpu.immdec.imm30_25[2] ;
 wire \u_cpu.cpu.immdec.imm30_25[3] ;
 wire \u_cpu.cpu.immdec.imm30_25[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[5] ;
 wire \u_cpu.cpu.immdec.imm31 ;
 wire \u_cpu.cpu.immdec.imm7 ;
 wire \u_cpu.cpu.mem_bytecnt[0] ;
 wire \u_cpu.cpu.mem_bytecnt[1] ;
 wire \u_cpu.cpu.mem_if.signbit ;
 wire \u_cpu.cpu.o_wdata0 ;
 wire \u_cpu.cpu.o_wdata1 ;
 wire \u_cpu.cpu.o_wen0 ;
 wire \u_cpu.cpu.o_wen1 ;
 wire \u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \u_cpu.cpu.state.ibus_cyc ;
 wire \u_cpu.cpu.state.init_done ;
 wire \u_cpu.cpu.state.o_cnt[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[0] ;
 wire \u_cpu.cpu.state.o_cnt_r[1] ;
 wire \u_cpu.cpu.state.o_cnt_r[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[3] ;
 wire \u_cpu.cpu.state.stage_two_req ;
 wire \u_cpu.raddr[0] ;
 wire \u_cpu.raddr[1] ;
 wire \u_cpu.rf_ram.memory[0][0] ;
 wire \u_cpu.rf_ram.memory[0][1] ;
 wire \u_cpu.rf_ram.memory[0][2] ;
 wire \u_cpu.rf_ram.memory[0][3] ;
 wire \u_cpu.rf_ram.memory[0][4] ;
 wire \u_cpu.rf_ram.memory[0][5] ;
 wire \u_cpu.rf_ram.memory[0][6] ;
 wire \u_cpu.rf_ram.memory[0][7] ;
 wire \u_cpu.rf_ram.memory[100][0] ;
 wire \u_cpu.rf_ram.memory[100][1] ;
 wire \u_cpu.rf_ram.memory[100][2] ;
 wire \u_cpu.rf_ram.memory[100][3] ;
 wire \u_cpu.rf_ram.memory[100][4] ;
 wire \u_cpu.rf_ram.memory[100][5] ;
 wire \u_cpu.rf_ram.memory[100][6] ;
 wire \u_cpu.rf_ram.memory[100][7] ;
 wire \u_cpu.rf_ram.memory[101][0] ;
 wire \u_cpu.rf_ram.memory[101][1] ;
 wire \u_cpu.rf_ram.memory[101][2] ;
 wire \u_cpu.rf_ram.memory[101][3] ;
 wire \u_cpu.rf_ram.memory[101][4] ;
 wire \u_cpu.rf_ram.memory[101][5] ;
 wire \u_cpu.rf_ram.memory[101][6] ;
 wire \u_cpu.rf_ram.memory[101][7] ;
 wire \u_cpu.rf_ram.memory[102][0] ;
 wire \u_cpu.rf_ram.memory[102][1] ;
 wire \u_cpu.rf_ram.memory[102][2] ;
 wire \u_cpu.rf_ram.memory[102][3] ;
 wire \u_cpu.rf_ram.memory[102][4] ;
 wire \u_cpu.rf_ram.memory[102][5] ;
 wire \u_cpu.rf_ram.memory[102][6] ;
 wire \u_cpu.rf_ram.memory[102][7] ;
 wire \u_cpu.rf_ram.memory[103][0] ;
 wire \u_cpu.rf_ram.memory[103][1] ;
 wire \u_cpu.rf_ram.memory[103][2] ;
 wire \u_cpu.rf_ram.memory[103][3] ;
 wire \u_cpu.rf_ram.memory[103][4] ;
 wire \u_cpu.rf_ram.memory[103][5] ;
 wire \u_cpu.rf_ram.memory[103][6] ;
 wire \u_cpu.rf_ram.memory[103][7] ;
 wire \u_cpu.rf_ram.memory[104][0] ;
 wire \u_cpu.rf_ram.memory[104][1] ;
 wire \u_cpu.rf_ram.memory[104][2] ;
 wire \u_cpu.rf_ram.memory[104][3] ;
 wire \u_cpu.rf_ram.memory[104][4] ;
 wire \u_cpu.rf_ram.memory[104][5] ;
 wire \u_cpu.rf_ram.memory[104][6] ;
 wire \u_cpu.rf_ram.memory[104][7] ;
 wire \u_cpu.rf_ram.memory[105][0] ;
 wire \u_cpu.rf_ram.memory[105][1] ;
 wire \u_cpu.rf_ram.memory[105][2] ;
 wire \u_cpu.rf_ram.memory[105][3] ;
 wire \u_cpu.rf_ram.memory[105][4] ;
 wire \u_cpu.rf_ram.memory[105][5] ;
 wire \u_cpu.rf_ram.memory[105][6] ;
 wire \u_cpu.rf_ram.memory[105][7] ;
 wire \u_cpu.rf_ram.memory[106][0] ;
 wire \u_cpu.rf_ram.memory[106][1] ;
 wire \u_cpu.rf_ram.memory[106][2] ;
 wire \u_cpu.rf_ram.memory[106][3] ;
 wire \u_cpu.rf_ram.memory[106][4] ;
 wire \u_cpu.rf_ram.memory[106][5] ;
 wire \u_cpu.rf_ram.memory[106][6] ;
 wire \u_cpu.rf_ram.memory[106][7] ;
 wire \u_cpu.rf_ram.memory[107][0] ;
 wire \u_cpu.rf_ram.memory[107][1] ;
 wire \u_cpu.rf_ram.memory[107][2] ;
 wire \u_cpu.rf_ram.memory[107][3] ;
 wire \u_cpu.rf_ram.memory[107][4] ;
 wire \u_cpu.rf_ram.memory[107][5] ;
 wire \u_cpu.rf_ram.memory[107][6] ;
 wire \u_cpu.rf_ram.memory[107][7] ;
 wire \u_cpu.rf_ram.memory[108][0] ;
 wire \u_cpu.rf_ram.memory[108][1] ;
 wire \u_cpu.rf_ram.memory[108][2] ;
 wire \u_cpu.rf_ram.memory[108][3] ;
 wire \u_cpu.rf_ram.memory[108][4] ;
 wire \u_cpu.rf_ram.memory[108][5] ;
 wire \u_cpu.rf_ram.memory[108][6] ;
 wire \u_cpu.rf_ram.memory[108][7] ;
 wire \u_cpu.rf_ram.memory[109][0] ;
 wire \u_cpu.rf_ram.memory[109][1] ;
 wire \u_cpu.rf_ram.memory[109][2] ;
 wire \u_cpu.rf_ram.memory[109][3] ;
 wire \u_cpu.rf_ram.memory[109][4] ;
 wire \u_cpu.rf_ram.memory[109][5] ;
 wire \u_cpu.rf_ram.memory[109][6] ;
 wire \u_cpu.rf_ram.memory[109][7] ;
 wire \u_cpu.rf_ram.memory[10][0] ;
 wire \u_cpu.rf_ram.memory[10][1] ;
 wire \u_cpu.rf_ram.memory[10][2] ;
 wire \u_cpu.rf_ram.memory[10][3] ;
 wire \u_cpu.rf_ram.memory[10][4] ;
 wire \u_cpu.rf_ram.memory[10][5] ;
 wire \u_cpu.rf_ram.memory[10][6] ;
 wire \u_cpu.rf_ram.memory[10][7] ;
 wire \u_cpu.rf_ram.memory[110][0] ;
 wire \u_cpu.rf_ram.memory[110][1] ;
 wire \u_cpu.rf_ram.memory[110][2] ;
 wire \u_cpu.rf_ram.memory[110][3] ;
 wire \u_cpu.rf_ram.memory[110][4] ;
 wire \u_cpu.rf_ram.memory[110][5] ;
 wire \u_cpu.rf_ram.memory[110][6] ;
 wire \u_cpu.rf_ram.memory[110][7] ;
 wire \u_cpu.rf_ram.memory[111][0] ;
 wire \u_cpu.rf_ram.memory[111][1] ;
 wire \u_cpu.rf_ram.memory[111][2] ;
 wire \u_cpu.rf_ram.memory[111][3] ;
 wire \u_cpu.rf_ram.memory[111][4] ;
 wire \u_cpu.rf_ram.memory[111][5] ;
 wire \u_cpu.rf_ram.memory[111][6] ;
 wire \u_cpu.rf_ram.memory[111][7] ;
 wire \u_cpu.rf_ram.memory[112][0] ;
 wire \u_cpu.rf_ram.memory[112][1] ;
 wire \u_cpu.rf_ram.memory[112][2] ;
 wire \u_cpu.rf_ram.memory[112][3] ;
 wire \u_cpu.rf_ram.memory[112][4] ;
 wire \u_cpu.rf_ram.memory[112][5] ;
 wire \u_cpu.rf_ram.memory[112][6] ;
 wire \u_cpu.rf_ram.memory[112][7] ;
 wire \u_cpu.rf_ram.memory[113][0] ;
 wire \u_cpu.rf_ram.memory[113][1] ;
 wire \u_cpu.rf_ram.memory[113][2] ;
 wire \u_cpu.rf_ram.memory[113][3] ;
 wire \u_cpu.rf_ram.memory[113][4] ;
 wire \u_cpu.rf_ram.memory[113][5] ;
 wire \u_cpu.rf_ram.memory[113][6] ;
 wire \u_cpu.rf_ram.memory[113][7] ;
 wire \u_cpu.rf_ram.memory[114][0] ;
 wire \u_cpu.rf_ram.memory[114][1] ;
 wire \u_cpu.rf_ram.memory[114][2] ;
 wire \u_cpu.rf_ram.memory[114][3] ;
 wire \u_cpu.rf_ram.memory[114][4] ;
 wire \u_cpu.rf_ram.memory[114][5] ;
 wire \u_cpu.rf_ram.memory[114][6] ;
 wire \u_cpu.rf_ram.memory[114][7] ;
 wire \u_cpu.rf_ram.memory[115][0] ;
 wire \u_cpu.rf_ram.memory[115][1] ;
 wire \u_cpu.rf_ram.memory[115][2] ;
 wire \u_cpu.rf_ram.memory[115][3] ;
 wire \u_cpu.rf_ram.memory[115][4] ;
 wire \u_cpu.rf_ram.memory[115][5] ;
 wire \u_cpu.rf_ram.memory[115][6] ;
 wire \u_cpu.rf_ram.memory[115][7] ;
 wire \u_cpu.rf_ram.memory[116][0] ;
 wire \u_cpu.rf_ram.memory[116][1] ;
 wire \u_cpu.rf_ram.memory[116][2] ;
 wire \u_cpu.rf_ram.memory[116][3] ;
 wire \u_cpu.rf_ram.memory[116][4] ;
 wire \u_cpu.rf_ram.memory[116][5] ;
 wire \u_cpu.rf_ram.memory[116][6] ;
 wire \u_cpu.rf_ram.memory[116][7] ;
 wire \u_cpu.rf_ram.memory[117][0] ;
 wire \u_cpu.rf_ram.memory[117][1] ;
 wire \u_cpu.rf_ram.memory[117][2] ;
 wire \u_cpu.rf_ram.memory[117][3] ;
 wire \u_cpu.rf_ram.memory[117][4] ;
 wire \u_cpu.rf_ram.memory[117][5] ;
 wire \u_cpu.rf_ram.memory[117][6] ;
 wire \u_cpu.rf_ram.memory[117][7] ;
 wire \u_cpu.rf_ram.memory[118][0] ;
 wire \u_cpu.rf_ram.memory[118][1] ;
 wire \u_cpu.rf_ram.memory[118][2] ;
 wire \u_cpu.rf_ram.memory[118][3] ;
 wire \u_cpu.rf_ram.memory[118][4] ;
 wire \u_cpu.rf_ram.memory[118][5] ;
 wire \u_cpu.rf_ram.memory[118][6] ;
 wire \u_cpu.rf_ram.memory[118][7] ;
 wire \u_cpu.rf_ram.memory[119][0] ;
 wire \u_cpu.rf_ram.memory[119][1] ;
 wire \u_cpu.rf_ram.memory[119][2] ;
 wire \u_cpu.rf_ram.memory[119][3] ;
 wire \u_cpu.rf_ram.memory[119][4] ;
 wire \u_cpu.rf_ram.memory[119][5] ;
 wire \u_cpu.rf_ram.memory[119][6] ;
 wire \u_cpu.rf_ram.memory[119][7] ;
 wire \u_cpu.rf_ram.memory[11][0] ;
 wire \u_cpu.rf_ram.memory[11][1] ;
 wire \u_cpu.rf_ram.memory[11][2] ;
 wire \u_cpu.rf_ram.memory[11][3] ;
 wire \u_cpu.rf_ram.memory[11][4] ;
 wire \u_cpu.rf_ram.memory[11][5] ;
 wire \u_cpu.rf_ram.memory[11][6] ;
 wire \u_cpu.rf_ram.memory[11][7] ;
 wire \u_cpu.rf_ram.memory[120][0] ;
 wire \u_cpu.rf_ram.memory[120][1] ;
 wire \u_cpu.rf_ram.memory[120][2] ;
 wire \u_cpu.rf_ram.memory[120][3] ;
 wire \u_cpu.rf_ram.memory[120][4] ;
 wire \u_cpu.rf_ram.memory[120][5] ;
 wire \u_cpu.rf_ram.memory[120][6] ;
 wire \u_cpu.rf_ram.memory[120][7] ;
 wire \u_cpu.rf_ram.memory[121][0] ;
 wire \u_cpu.rf_ram.memory[121][1] ;
 wire \u_cpu.rf_ram.memory[121][2] ;
 wire \u_cpu.rf_ram.memory[121][3] ;
 wire \u_cpu.rf_ram.memory[121][4] ;
 wire \u_cpu.rf_ram.memory[121][5] ;
 wire \u_cpu.rf_ram.memory[121][6] ;
 wire \u_cpu.rf_ram.memory[121][7] ;
 wire \u_cpu.rf_ram.memory[122][0] ;
 wire \u_cpu.rf_ram.memory[122][1] ;
 wire \u_cpu.rf_ram.memory[122][2] ;
 wire \u_cpu.rf_ram.memory[122][3] ;
 wire \u_cpu.rf_ram.memory[122][4] ;
 wire \u_cpu.rf_ram.memory[122][5] ;
 wire \u_cpu.rf_ram.memory[122][6] ;
 wire \u_cpu.rf_ram.memory[122][7] ;
 wire \u_cpu.rf_ram.memory[123][0] ;
 wire \u_cpu.rf_ram.memory[123][1] ;
 wire \u_cpu.rf_ram.memory[123][2] ;
 wire \u_cpu.rf_ram.memory[123][3] ;
 wire \u_cpu.rf_ram.memory[123][4] ;
 wire \u_cpu.rf_ram.memory[123][5] ;
 wire \u_cpu.rf_ram.memory[123][6] ;
 wire \u_cpu.rf_ram.memory[123][7] ;
 wire \u_cpu.rf_ram.memory[124][0] ;
 wire \u_cpu.rf_ram.memory[124][1] ;
 wire \u_cpu.rf_ram.memory[124][2] ;
 wire \u_cpu.rf_ram.memory[124][3] ;
 wire \u_cpu.rf_ram.memory[124][4] ;
 wire \u_cpu.rf_ram.memory[124][5] ;
 wire \u_cpu.rf_ram.memory[124][6] ;
 wire \u_cpu.rf_ram.memory[124][7] ;
 wire \u_cpu.rf_ram.memory[125][0] ;
 wire \u_cpu.rf_ram.memory[125][1] ;
 wire \u_cpu.rf_ram.memory[125][2] ;
 wire \u_cpu.rf_ram.memory[125][3] ;
 wire \u_cpu.rf_ram.memory[125][4] ;
 wire \u_cpu.rf_ram.memory[125][5] ;
 wire \u_cpu.rf_ram.memory[125][6] ;
 wire \u_cpu.rf_ram.memory[125][7] ;
 wire \u_cpu.rf_ram.memory[126][0] ;
 wire \u_cpu.rf_ram.memory[126][1] ;
 wire \u_cpu.rf_ram.memory[126][2] ;
 wire \u_cpu.rf_ram.memory[126][3] ;
 wire \u_cpu.rf_ram.memory[126][4] ;
 wire \u_cpu.rf_ram.memory[126][5] ;
 wire \u_cpu.rf_ram.memory[126][6] ;
 wire \u_cpu.rf_ram.memory[126][7] ;
 wire \u_cpu.rf_ram.memory[127][0] ;
 wire \u_cpu.rf_ram.memory[127][1] ;
 wire \u_cpu.rf_ram.memory[127][2] ;
 wire \u_cpu.rf_ram.memory[127][3] ;
 wire \u_cpu.rf_ram.memory[127][4] ;
 wire \u_cpu.rf_ram.memory[127][5] ;
 wire \u_cpu.rf_ram.memory[127][6] ;
 wire \u_cpu.rf_ram.memory[127][7] ;
 wire \u_cpu.rf_ram.memory[128][0] ;
 wire \u_cpu.rf_ram.memory[128][1] ;
 wire \u_cpu.rf_ram.memory[128][2] ;
 wire \u_cpu.rf_ram.memory[128][3] ;
 wire \u_cpu.rf_ram.memory[128][4] ;
 wire \u_cpu.rf_ram.memory[128][5] ;
 wire \u_cpu.rf_ram.memory[128][6] ;
 wire \u_cpu.rf_ram.memory[128][7] ;
 wire \u_cpu.rf_ram.memory[129][0] ;
 wire \u_cpu.rf_ram.memory[129][1] ;
 wire \u_cpu.rf_ram.memory[129][2] ;
 wire \u_cpu.rf_ram.memory[129][3] ;
 wire \u_cpu.rf_ram.memory[129][4] ;
 wire \u_cpu.rf_ram.memory[129][5] ;
 wire \u_cpu.rf_ram.memory[129][6] ;
 wire \u_cpu.rf_ram.memory[129][7] ;
 wire \u_cpu.rf_ram.memory[12][0] ;
 wire \u_cpu.rf_ram.memory[12][1] ;
 wire \u_cpu.rf_ram.memory[12][2] ;
 wire \u_cpu.rf_ram.memory[12][3] ;
 wire \u_cpu.rf_ram.memory[12][4] ;
 wire \u_cpu.rf_ram.memory[12][5] ;
 wire \u_cpu.rf_ram.memory[12][6] ;
 wire \u_cpu.rf_ram.memory[12][7] ;
 wire \u_cpu.rf_ram.memory[130][0] ;
 wire \u_cpu.rf_ram.memory[130][1] ;
 wire \u_cpu.rf_ram.memory[130][2] ;
 wire \u_cpu.rf_ram.memory[130][3] ;
 wire \u_cpu.rf_ram.memory[130][4] ;
 wire \u_cpu.rf_ram.memory[130][5] ;
 wire \u_cpu.rf_ram.memory[130][6] ;
 wire \u_cpu.rf_ram.memory[130][7] ;
 wire \u_cpu.rf_ram.memory[131][0] ;
 wire \u_cpu.rf_ram.memory[131][1] ;
 wire \u_cpu.rf_ram.memory[131][2] ;
 wire \u_cpu.rf_ram.memory[131][3] ;
 wire \u_cpu.rf_ram.memory[131][4] ;
 wire \u_cpu.rf_ram.memory[131][5] ;
 wire \u_cpu.rf_ram.memory[131][6] ;
 wire \u_cpu.rf_ram.memory[131][7] ;
 wire \u_cpu.rf_ram.memory[132][0] ;
 wire \u_cpu.rf_ram.memory[132][1] ;
 wire \u_cpu.rf_ram.memory[132][2] ;
 wire \u_cpu.rf_ram.memory[132][3] ;
 wire \u_cpu.rf_ram.memory[132][4] ;
 wire \u_cpu.rf_ram.memory[132][5] ;
 wire \u_cpu.rf_ram.memory[132][6] ;
 wire \u_cpu.rf_ram.memory[132][7] ;
 wire \u_cpu.rf_ram.memory[133][0] ;
 wire \u_cpu.rf_ram.memory[133][1] ;
 wire \u_cpu.rf_ram.memory[133][2] ;
 wire \u_cpu.rf_ram.memory[133][3] ;
 wire \u_cpu.rf_ram.memory[133][4] ;
 wire \u_cpu.rf_ram.memory[133][5] ;
 wire \u_cpu.rf_ram.memory[133][6] ;
 wire \u_cpu.rf_ram.memory[133][7] ;
 wire \u_cpu.rf_ram.memory[134][0] ;
 wire \u_cpu.rf_ram.memory[134][1] ;
 wire \u_cpu.rf_ram.memory[134][2] ;
 wire \u_cpu.rf_ram.memory[134][3] ;
 wire \u_cpu.rf_ram.memory[134][4] ;
 wire \u_cpu.rf_ram.memory[134][5] ;
 wire \u_cpu.rf_ram.memory[134][6] ;
 wire \u_cpu.rf_ram.memory[134][7] ;
 wire \u_cpu.rf_ram.memory[135][0] ;
 wire \u_cpu.rf_ram.memory[135][1] ;
 wire \u_cpu.rf_ram.memory[135][2] ;
 wire \u_cpu.rf_ram.memory[135][3] ;
 wire \u_cpu.rf_ram.memory[135][4] ;
 wire \u_cpu.rf_ram.memory[135][5] ;
 wire \u_cpu.rf_ram.memory[135][6] ;
 wire \u_cpu.rf_ram.memory[135][7] ;
 wire \u_cpu.rf_ram.memory[136][0] ;
 wire \u_cpu.rf_ram.memory[136][1] ;
 wire \u_cpu.rf_ram.memory[136][2] ;
 wire \u_cpu.rf_ram.memory[136][3] ;
 wire \u_cpu.rf_ram.memory[136][4] ;
 wire \u_cpu.rf_ram.memory[136][5] ;
 wire \u_cpu.rf_ram.memory[136][6] ;
 wire \u_cpu.rf_ram.memory[136][7] ;
 wire \u_cpu.rf_ram.memory[137][0] ;
 wire \u_cpu.rf_ram.memory[137][1] ;
 wire \u_cpu.rf_ram.memory[137][2] ;
 wire \u_cpu.rf_ram.memory[137][3] ;
 wire \u_cpu.rf_ram.memory[137][4] ;
 wire \u_cpu.rf_ram.memory[137][5] ;
 wire \u_cpu.rf_ram.memory[137][6] ;
 wire \u_cpu.rf_ram.memory[137][7] ;
 wire \u_cpu.rf_ram.memory[138][0] ;
 wire \u_cpu.rf_ram.memory[138][1] ;
 wire \u_cpu.rf_ram.memory[138][2] ;
 wire \u_cpu.rf_ram.memory[138][3] ;
 wire \u_cpu.rf_ram.memory[138][4] ;
 wire \u_cpu.rf_ram.memory[138][5] ;
 wire \u_cpu.rf_ram.memory[138][6] ;
 wire \u_cpu.rf_ram.memory[138][7] ;
 wire \u_cpu.rf_ram.memory[139][0] ;
 wire \u_cpu.rf_ram.memory[139][1] ;
 wire \u_cpu.rf_ram.memory[139][2] ;
 wire \u_cpu.rf_ram.memory[139][3] ;
 wire \u_cpu.rf_ram.memory[139][4] ;
 wire \u_cpu.rf_ram.memory[139][5] ;
 wire \u_cpu.rf_ram.memory[139][6] ;
 wire \u_cpu.rf_ram.memory[139][7] ;
 wire \u_cpu.rf_ram.memory[13][0] ;
 wire \u_cpu.rf_ram.memory[13][1] ;
 wire \u_cpu.rf_ram.memory[13][2] ;
 wire \u_cpu.rf_ram.memory[13][3] ;
 wire \u_cpu.rf_ram.memory[13][4] ;
 wire \u_cpu.rf_ram.memory[13][5] ;
 wire \u_cpu.rf_ram.memory[13][6] ;
 wire \u_cpu.rf_ram.memory[13][7] ;
 wire \u_cpu.rf_ram.memory[140][0] ;
 wire \u_cpu.rf_ram.memory[140][1] ;
 wire \u_cpu.rf_ram.memory[140][2] ;
 wire \u_cpu.rf_ram.memory[140][3] ;
 wire \u_cpu.rf_ram.memory[140][4] ;
 wire \u_cpu.rf_ram.memory[140][5] ;
 wire \u_cpu.rf_ram.memory[140][6] ;
 wire \u_cpu.rf_ram.memory[140][7] ;
 wire \u_cpu.rf_ram.memory[141][0] ;
 wire \u_cpu.rf_ram.memory[141][1] ;
 wire \u_cpu.rf_ram.memory[141][2] ;
 wire \u_cpu.rf_ram.memory[141][3] ;
 wire \u_cpu.rf_ram.memory[141][4] ;
 wire \u_cpu.rf_ram.memory[141][5] ;
 wire \u_cpu.rf_ram.memory[141][6] ;
 wire \u_cpu.rf_ram.memory[141][7] ;
 wire \u_cpu.rf_ram.memory[142][0] ;
 wire \u_cpu.rf_ram.memory[142][1] ;
 wire \u_cpu.rf_ram.memory[142][2] ;
 wire \u_cpu.rf_ram.memory[142][3] ;
 wire \u_cpu.rf_ram.memory[142][4] ;
 wire \u_cpu.rf_ram.memory[142][5] ;
 wire \u_cpu.rf_ram.memory[142][6] ;
 wire \u_cpu.rf_ram.memory[142][7] ;
 wire \u_cpu.rf_ram.memory[143][0] ;
 wire \u_cpu.rf_ram.memory[143][1] ;
 wire \u_cpu.rf_ram.memory[143][2] ;
 wire \u_cpu.rf_ram.memory[143][3] ;
 wire \u_cpu.rf_ram.memory[143][4] ;
 wire \u_cpu.rf_ram.memory[143][5] ;
 wire \u_cpu.rf_ram.memory[143][6] ;
 wire \u_cpu.rf_ram.memory[143][7] ;
 wire \u_cpu.rf_ram.memory[14][0] ;
 wire \u_cpu.rf_ram.memory[14][1] ;
 wire \u_cpu.rf_ram.memory[14][2] ;
 wire \u_cpu.rf_ram.memory[14][3] ;
 wire \u_cpu.rf_ram.memory[14][4] ;
 wire \u_cpu.rf_ram.memory[14][5] ;
 wire \u_cpu.rf_ram.memory[14][6] ;
 wire \u_cpu.rf_ram.memory[14][7] ;
 wire \u_cpu.rf_ram.memory[15][0] ;
 wire \u_cpu.rf_ram.memory[15][1] ;
 wire \u_cpu.rf_ram.memory[15][2] ;
 wire \u_cpu.rf_ram.memory[15][3] ;
 wire \u_cpu.rf_ram.memory[15][4] ;
 wire \u_cpu.rf_ram.memory[15][5] ;
 wire \u_cpu.rf_ram.memory[15][6] ;
 wire \u_cpu.rf_ram.memory[15][7] ;
 wire \u_cpu.rf_ram.memory[16][0] ;
 wire \u_cpu.rf_ram.memory[16][1] ;
 wire \u_cpu.rf_ram.memory[16][2] ;
 wire \u_cpu.rf_ram.memory[16][3] ;
 wire \u_cpu.rf_ram.memory[16][4] ;
 wire \u_cpu.rf_ram.memory[16][5] ;
 wire \u_cpu.rf_ram.memory[16][6] ;
 wire \u_cpu.rf_ram.memory[16][7] ;
 wire \u_cpu.rf_ram.memory[17][0] ;
 wire \u_cpu.rf_ram.memory[17][1] ;
 wire \u_cpu.rf_ram.memory[17][2] ;
 wire \u_cpu.rf_ram.memory[17][3] ;
 wire \u_cpu.rf_ram.memory[17][4] ;
 wire \u_cpu.rf_ram.memory[17][5] ;
 wire \u_cpu.rf_ram.memory[17][6] ;
 wire \u_cpu.rf_ram.memory[17][7] ;
 wire \u_cpu.rf_ram.memory[18][0] ;
 wire \u_cpu.rf_ram.memory[18][1] ;
 wire \u_cpu.rf_ram.memory[18][2] ;
 wire \u_cpu.rf_ram.memory[18][3] ;
 wire \u_cpu.rf_ram.memory[18][4] ;
 wire \u_cpu.rf_ram.memory[18][5] ;
 wire \u_cpu.rf_ram.memory[18][6] ;
 wire \u_cpu.rf_ram.memory[18][7] ;
 wire \u_cpu.rf_ram.memory[19][0] ;
 wire \u_cpu.rf_ram.memory[19][1] ;
 wire \u_cpu.rf_ram.memory[19][2] ;
 wire \u_cpu.rf_ram.memory[19][3] ;
 wire \u_cpu.rf_ram.memory[19][4] ;
 wire \u_cpu.rf_ram.memory[19][5] ;
 wire \u_cpu.rf_ram.memory[19][6] ;
 wire \u_cpu.rf_ram.memory[19][7] ;
 wire \u_cpu.rf_ram.memory[1][0] ;
 wire \u_cpu.rf_ram.memory[1][1] ;
 wire \u_cpu.rf_ram.memory[1][2] ;
 wire \u_cpu.rf_ram.memory[1][3] ;
 wire \u_cpu.rf_ram.memory[1][4] ;
 wire \u_cpu.rf_ram.memory[1][5] ;
 wire \u_cpu.rf_ram.memory[1][6] ;
 wire \u_cpu.rf_ram.memory[1][7] ;
 wire \u_cpu.rf_ram.memory[20][0] ;
 wire \u_cpu.rf_ram.memory[20][1] ;
 wire \u_cpu.rf_ram.memory[20][2] ;
 wire \u_cpu.rf_ram.memory[20][3] ;
 wire \u_cpu.rf_ram.memory[20][4] ;
 wire \u_cpu.rf_ram.memory[20][5] ;
 wire \u_cpu.rf_ram.memory[20][6] ;
 wire \u_cpu.rf_ram.memory[20][7] ;
 wire \u_cpu.rf_ram.memory[21][0] ;
 wire \u_cpu.rf_ram.memory[21][1] ;
 wire \u_cpu.rf_ram.memory[21][2] ;
 wire \u_cpu.rf_ram.memory[21][3] ;
 wire \u_cpu.rf_ram.memory[21][4] ;
 wire \u_cpu.rf_ram.memory[21][5] ;
 wire \u_cpu.rf_ram.memory[21][6] ;
 wire \u_cpu.rf_ram.memory[21][7] ;
 wire \u_cpu.rf_ram.memory[22][0] ;
 wire \u_cpu.rf_ram.memory[22][1] ;
 wire \u_cpu.rf_ram.memory[22][2] ;
 wire \u_cpu.rf_ram.memory[22][3] ;
 wire \u_cpu.rf_ram.memory[22][4] ;
 wire \u_cpu.rf_ram.memory[22][5] ;
 wire \u_cpu.rf_ram.memory[22][6] ;
 wire \u_cpu.rf_ram.memory[22][7] ;
 wire \u_cpu.rf_ram.memory[23][0] ;
 wire \u_cpu.rf_ram.memory[23][1] ;
 wire \u_cpu.rf_ram.memory[23][2] ;
 wire \u_cpu.rf_ram.memory[23][3] ;
 wire \u_cpu.rf_ram.memory[23][4] ;
 wire \u_cpu.rf_ram.memory[23][5] ;
 wire \u_cpu.rf_ram.memory[23][6] ;
 wire \u_cpu.rf_ram.memory[23][7] ;
 wire \u_cpu.rf_ram.memory[24][0] ;
 wire \u_cpu.rf_ram.memory[24][1] ;
 wire \u_cpu.rf_ram.memory[24][2] ;
 wire \u_cpu.rf_ram.memory[24][3] ;
 wire \u_cpu.rf_ram.memory[24][4] ;
 wire \u_cpu.rf_ram.memory[24][5] ;
 wire \u_cpu.rf_ram.memory[24][6] ;
 wire \u_cpu.rf_ram.memory[24][7] ;
 wire \u_cpu.rf_ram.memory[25][0] ;
 wire \u_cpu.rf_ram.memory[25][1] ;
 wire \u_cpu.rf_ram.memory[25][2] ;
 wire \u_cpu.rf_ram.memory[25][3] ;
 wire \u_cpu.rf_ram.memory[25][4] ;
 wire \u_cpu.rf_ram.memory[25][5] ;
 wire \u_cpu.rf_ram.memory[25][6] ;
 wire \u_cpu.rf_ram.memory[25][7] ;
 wire \u_cpu.rf_ram.memory[26][0] ;
 wire \u_cpu.rf_ram.memory[26][1] ;
 wire \u_cpu.rf_ram.memory[26][2] ;
 wire \u_cpu.rf_ram.memory[26][3] ;
 wire \u_cpu.rf_ram.memory[26][4] ;
 wire \u_cpu.rf_ram.memory[26][5] ;
 wire \u_cpu.rf_ram.memory[26][6] ;
 wire \u_cpu.rf_ram.memory[26][7] ;
 wire \u_cpu.rf_ram.memory[27][0] ;
 wire \u_cpu.rf_ram.memory[27][1] ;
 wire \u_cpu.rf_ram.memory[27][2] ;
 wire \u_cpu.rf_ram.memory[27][3] ;
 wire \u_cpu.rf_ram.memory[27][4] ;
 wire \u_cpu.rf_ram.memory[27][5] ;
 wire \u_cpu.rf_ram.memory[27][6] ;
 wire \u_cpu.rf_ram.memory[27][7] ;
 wire \u_cpu.rf_ram.memory[28][0] ;
 wire \u_cpu.rf_ram.memory[28][1] ;
 wire \u_cpu.rf_ram.memory[28][2] ;
 wire \u_cpu.rf_ram.memory[28][3] ;
 wire \u_cpu.rf_ram.memory[28][4] ;
 wire \u_cpu.rf_ram.memory[28][5] ;
 wire \u_cpu.rf_ram.memory[28][6] ;
 wire \u_cpu.rf_ram.memory[28][7] ;
 wire \u_cpu.rf_ram.memory[29][0] ;
 wire \u_cpu.rf_ram.memory[29][1] ;
 wire \u_cpu.rf_ram.memory[29][2] ;
 wire \u_cpu.rf_ram.memory[29][3] ;
 wire \u_cpu.rf_ram.memory[29][4] ;
 wire \u_cpu.rf_ram.memory[29][5] ;
 wire \u_cpu.rf_ram.memory[29][6] ;
 wire \u_cpu.rf_ram.memory[29][7] ;
 wire \u_cpu.rf_ram.memory[2][0] ;
 wire \u_cpu.rf_ram.memory[2][1] ;
 wire \u_cpu.rf_ram.memory[2][2] ;
 wire \u_cpu.rf_ram.memory[2][3] ;
 wire \u_cpu.rf_ram.memory[2][4] ;
 wire \u_cpu.rf_ram.memory[2][5] ;
 wire \u_cpu.rf_ram.memory[2][6] ;
 wire \u_cpu.rf_ram.memory[2][7] ;
 wire \u_cpu.rf_ram.memory[30][0] ;
 wire \u_cpu.rf_ram.memory[30][1] ;
 wire \u_cpu.rf_ram.memory[30][2] ;
 wire \u_cpu.rf_ram.memory[30][3] ;
 wire \u_cpu.rf_ram.memory[30][4] ;
 wire \u_cpu.rf_ram.memory[30][5] ;
 wire \u_cpu.rf_ram.memory[30][6] ;
 wire \u_cpu.rf_ram.memory[30][7] ;
 wire \u_cpu.rf_ram.memory[31][0] ;
 wire \u_cpu.rf_ram.memory[31][1] ;
 wire \u_cpu.rf_ram.memory[31][2] ;
 wire \u_cpu.rf_ram.memory[31][3] ;
 wire \u_cpu.rf_ram.memory[31][4] ;
 wire \u_cpu.rf_ram.memory[31][5] ;
 wire \u_cpu.rf_ram.memory[31][6] ;
 wire \u_cpu.rf_ram.memory[31][7] ;
 wire \u_cpu.rf_ram.memory[32][0] ;
 wire \u_cpu.rf_ram.memory[32][1] ;
 wire \u_cpu.rf_ram.memory[32][2] ;
 wire \u_cpu.rf_ram.memory[32][3] ;
 wire \u_cpu.rf_ram.memory[32][4] ;
 wire \u_cpu.rf_ram.memory[32][5] ;
 wire \u_cpu.rf_ram.memory[32][6] ;
 wire \u_cpu.rf_ram.memory[32][7] ;
 wire \u_cpu.rf_ram.memory[33][0] ;
 wire \u_cpu.rf_ram.memory[33][1] ;
 wire \u_cpu.rf_ram.memory[33][2] ;
 wire \u_cpu.rf_ram.memory[33][3] ;
 wire \u_cpu.rf_ram.memory[33][4] ;
 wire \u_cpu.rf_ram.memory[33][5] ;
 wire \u_cpu.rf_ram.memory[33][6] ;
 wire \u_cpu.rf_ram.memory[33][7] ;
 wire \u_cpu.rf_ram.memory[34][0] ;
 wire \u_cpu.rf_ram.memory[34][1] ;
 wire \u_cpu.rf_ram.memory[34][2] ;
 wire \u_cpu.rf_ram.memory[34][3] ;
 wire \u_cpu.rf_ram.memory[34][4] ;
 wire \u_cpu.rf_ram.memory[34][5] ;
 wire \u_cpu.rf_ram.memory[34][6] ;
 wire \u_cpu.rf_ram.memory[34][7] ;
 wire \u_cpu.rf_ram.memory[35][0] ;
 wire \u_cpu.rf_ram.memory[35][1] ;
 wire \u_cpu.rf_ram.memory[35][2] ;
 wire \u_cpu.rf_ram.memory[35][3] ;
 wire \u_cpu.rf_ram.memory[35][4] ;
 wire \u_cpu.rf_ram.memory[35][5] ;
 wire \u_cpu.rf_ram.memory[35][6] ;
 wire \u_cpu.rf_ram.memory[35][7] ;
 wire \u_cpu.rf_ram.memory[36][0] ;
 wire \u_cpu.rf_ram.memory[36][1] ;
 wire \u_cpu.rf_ram.memory[36][2] ;
 wire \u_cpu.rf_ram.memory[36][3] ;
 wire \u_cpu.rf_ram.memory[36][4] ;
 wire \u_cpu.rf_ram.memory[36][5] ;
 wire \u_cpu.rf_ram.memory[36][6] ;
 wire \u_cpu.rf_ram.memory[36][7] ;
 wire \u_cpu.rf_ram.memory[37][0] ;
 wire \u_cpu.rf_ram.memory[37][1] ;
 wire \u_cpu.rf_ram.memory[37][2] ;
 wire \u_cpu.rf_ram.memory[37][3] ;
 wire \u_cpu.rf_ram.memory[37][4] ;
 wire \u_cpu.rf_ram.memory[37][5] ;
 wire \u_cpu.rf_ram.memory[37][6] ;
 wire \u_cpu.rf_ram.memory[37][7] ;
 wire \u_cpu.rf_ram.memory[38][0] ;
 wire \u_cpu.rf_ram.memory[38][1] ;
 wire \u_cpu.rf_ram.memory[38][2] ;
 wire \u_cpu.rf_ram.memory[38][3] ;
 wire \u_cpu.rf_ram.memory[38][4] ;
 wire \u_cpu.rf_ram.memory[38][5] ;
 wire \u_cpu.rf_ram.memory[38][6] ;
 wire \u_cpu.rf_ram.memory[38][7] ;
 wire \u_cpu.rf_ram.memory[39][0] ;
 wire \u_cpu.rf_ram.memory[39][1] ;
 wire \u_cpu.rf_ram.memory[39][2] ;
 wire \u_cpu.rf_ram.memory[39][3] ;
 wire \u_cpu.rf_ram.memory[39][4] ;
 wire \u_cpu.rf_ram.memory[39][5] ;
 wire \u_cpu.rf_ram.memory[39][6] ;
 wire \u_cpu.rf_ram.memory[39][7] ;
 wire \u_cpu.rf_ram.memory[3][0] ;
 wire \u_cpu.rf_ram.memory[3][1] ;
 wire \u_cpu.rf_ram.memory[3][2] ;
 wire \u_cpu.rf_ram.memory[3][3] ;
 wire \u_cpu.rf_ram.memory[3][4] ;
 wire \u_cpu.rf_ram.memory[3][5] ;
 wire \u_cpu.rf_ram.memory[3][6] ;
 wire \u_cpu.rf_ram.memory[3][7] ;
 wire \u_cpu.rf_ram.memory[40][0] ;
 wire \u_cpu.rf_ram.memory[40][1] ;
 wire \u_cpu.rf_ram.memory[40][2] ;
 wire \u_cpu.rf_ram.memory[40][3] ;
 wire \u_cpu.rf_ram.memory[40][4] ;
 wire \u_cpu.rf_ram.memory[40][5] ;
 wire \u_cpu.rf_ram.memory[40][6] ;
 wire \u_cpu.rf_ram.memory[40][7] ;
 wire \u_cpu.rf_ram.memory[41][0] ;
 wire \u_cpu.rf_ram.memory[41][1] ;
 wire \u_cpu.rf_ram.memory[41][2] ;
 wire \u_cpu.rf_ram.memory[41][3] ;
 wire \u_cpu.rf_ram.memory[41][4] ;
 wire \u_cpu.rf_ram.memory[41][5] ;
 wire \u_cpu.rf_ram.memory[41][6] ;
 wire \u_cpu.rf_ram.memory[41][7] ;
 wire \u_cpu.rf_ram.memory[42][0] ;
 wire \u_cpu.rf_ram.memory[42][1] ;
 wire \u_cpu.rf_ram.memory[42][2] ;
 wire \u_cpu.rf_ram.memory[42][3] ;
 wire \u_cpu.rf_ram.memory[42][4] ;
 wire \u_cpu.rf_ram.memory[42][5] ;
 wire \u_cpu.rf_ram.memory[42][6] ;
 wire \u_cpu.rf_ram.memory[42][7] ;
 wire \u_cpu.rf_ram.memory[43][0] ;
 wire \u_cpu.rf_ram.memory[43][1] ;
 wire \u_cpu.rf_ram.memory[43][2] ;
 wire \u_cpu.rf_ram.memory[43][3] ;
 wire \u_cpu.rf_ram.memory[43][4] ;
 wire \u_cpu.rf_ram.memory[43][5] ;
 wire \u_cpu.rf_ram.memory[43][6] ;
 wire \u_cpu.rf_ram.memory[43][7] ;
 wire \u_cpu.rf_ram.memory[44][0] ;
 wire \u_cpu.rf_ram.memory[44][1] ;
 wire \u_cpu.rf_ram.memory[44][2] ;
 wire \u_cpu.rf_ram.memory[44][3] ;
 wire \u_cpu.rf_ram.memory[44][4] ;
 wire \u_cpu.rf_ram.memory[44][5] ;
 wire \u_cpu.rf_ram.memory[44][6] ;
 wire \u_cpu.rf_ram.memory[44][7] ;
 wire \u_cpu.rf_ram.memory[45][0] ;
 wire \u_cpu.rf_ram.memory[45][1] ;
 wire \u_cpu.rf_ram.memory[45][2] ;
 wire \u_cpu.rf_ram.memory[45][3] ;
 wire \u_cpu.rf_ram.memory[45][4] ;
 wire \u_cpu.rf_ram.memory[45][5] ;
 wire \u_cpu.rf_ram.memory[45][6] ;
 wire \u_cpu.rf_ram.memory[45][7] ;
 wire \u_cpu.rf_ram.memory[46][0] ;
 wire \u_cpu.rf_ram.memory[46][1] ;
 wire \u_cpu.rf_ram.memory[46][2] ;
 wire \u_cpu.rf_ram.memory[46][3] ;
 wire \u_cpu.rf_ram.memory[46][4] ;
 wire \u_cpu.rf_ram.memory[46][5] ;
 wire \u_cpu.rf_ram.memory[46][6] ;
 wire \u_cpu.rf_ram.memory[46][7] ;
 wire \u_cpu.rf_ram.memory[47][0] ;
 wire \u_cpu.rf_ram.memory[47][1] ;
 wire \u_cpu.rf_ram.memory[47][2] ;
 wire \u_cpu.rf_ram.memory[47][3] ;
 wire \u_cpu.rf_ram.memory[47][4] ;
 wire \u_cpu.rf_ram.memory[47][5] ;
 wire \u_cpu.rf_ram.memory[47][6] ;
 wire \u_cpu.rf_ram.memory[47][7] ;
 wire \u_cpu.rf_ram.memory[48][0] ;
 wire \u_cpu.rf_ram.memory[48][1] ;
 wire \u_cpu.rf_ram.memory[48][2] ;
 wire \u_cpu.rf_ram.memory[48][3] ;
 wire \u_cpu.rf_ram.memory[48][4] ;
 wire \u_cpu.rf_ram.memory[48][5] ;
 wire \u_cpu.rf_ram.memory[48][6] ;
 wire \u_cpu.rf_ram.memory[48][7] ;
 wire \u_cpu.rf_ram.memory[49][0] ;
 wire \u_cpu.rf_ram.memory[49][1] ;
 wire \u_cpu.rf_ram.memory[49][2] ;
 wire \u_cpu.rf_ram.memory[49][3] ;
 wire \u_cpu.rf_ram.memory[49][4] ;
 wire \u_cpu.rf_ram.memory[49][5] ;
 wire \u_cpu.rf_ram.memory[49][6] ;
 wire \u_cpu.rf_ram.memory[49][7] ;
 wire \u_cpu.rf_ram.memory[4][0] ;
 wire \u_cpu.rf_ram.memory[4][1] ;
 wire \u_cpu.rf_ram.memory[4][2] ;
 wire \u_cpu.rf_ram.memory[4][3] ;
 wire \u_cpu.rf_ram.memory[4][4] ;
 wire \u_cpu.rf_ram.memory[4][5] ;
 wire \u_cpu.rf_ram.memory[4][6] ;
 wire \u_cpu.rf_ram.memory[4][7] ;
 wire \u_cpu.rf_ram.memory[50][0] ;
 wire \u_cpu.rf_ram.memory[50][1] ;
 wire \u_cpu.rf_ram.memory[50][2] ;
 wire \u_cpu.rf_ram.memory[50][3] ;
 wire \u_cpu.rf_ram.memory[50][4] ;
 wire \u_cpu.rf_ram.memory[50][5] ;
 wire \u_cpu.rf_ram.memory[50][6] ;
 wire \u_cpu.rf_ram.memory[50][7] ;
 wire \u_cpu.rf_ram.memory[51][0] ;
 wire \u_cpu.rf_ram.memory[51][1] ;
 wire \u_cpu.rf_ram.memory[51][2] ;
 wire \u_cpu.rf_ram.memory[51][3] ;
 wire \u_cpu.rf_ram.memory[51][4] ;
 wire \u_cpu.rf_ram.memory[51][5] ;
 wire \u_cpu.rf_ram.memory[51][6] ;
 wire \u_cpu.rf_ram.memory[51][7] ;
 wire \u_cpu.rf_ram.memory[52][0] ;
 wire \u_cpu.rf_ram.memory[52][1] ;
 wire \u_cpu.rf_ram.memory[52][2] ;
 wire \u_cpu.rf_ram.memory[52][3] ;
 wire \u_cpu.rf_ram.memory[52][4] ;
 wire \u_cpu.rf_ram.memory[52][5] ;
 wire \u_cpu.rf_ram.memory[52][6] ;
 wire \u_cpu.rf_ram.memory[52][7] ;
 wire \u_cpu.rf_ram.memory[53][0] ;
 wire \u_cpu.rf_ram.memory[53][1] ;
 wire \u_cpu.rf_ram.memory[53][2] ;
 wire \u_cpu.rf_ram.memory[53][3] ;
 wire \u_cpu.rf_ram.memory[53][4] ;
 wire \u_cpu.rf_ram.memory[53][5] ;
 wire \u_cpu.rf_ram.memory[53][6] ;
 wire \u_cpu.rf_ram.memory[53][7] ;
 wire \u_cpu.rf_ram.memory[54][0] ;
 wire \u_cpu.rf_ram.memory[54][1] ;
 wire \u_cpu.rf_ram.memory[54][2] ;
 wire \u_cpu.rf_ram.memory[54][3] ;
 wire \u_cpu.rf_ram.memory[54][4] ;
 wire \u_cpu.rf_ram.memory[54][5] ;
 wire \u_cpu.rf_ram.memory[54][6] ;
 wire \u_cpu.rf_ram.memory[54][7] ;
 wire \u_cpu.rf_ram.memory[55][0] ;
 wire \u_cpu.rf_ram.memory[55][1] ;
 wire \u_cpu.rf_ram.memory[55][2] ;
 wire \u_cpu.rf_ram.memory[55][3] ;
 wire \u_cpu.rf_ram.memory[55][4] ;
 wire \u_cpu.rf_ram.memory[55][5] ;
 wire \u_cpu.rf_ram.memory[55][6] ;
 wire \u_cpu.rf_ram.memory[55][7] ;
 wire \u_cpu.rf_ram.memory[56][0] ;
 wire \u_cpu.rf_ram.memory[56][1] ;
 wire \u_cpu.rf_ram.memory[56][2] ;
 wire \u_cpu.rf_ram.memory[56][3] ;
 wire \u_cpu.rf_ram.memory[56][4] ;
 wire \u_cpu.rf_ram.memory[56][5] ;
 wire \u_cpu.rf_ram.memory[56][6] ;
 wire \u_cpu.rf_ram.memory[56][7] ;
 wire \u_cpu.rf_ram.memory[57][0] ;
 wire \u_cpu.rf_ram.memory[57][1] ;
 wire \u_cpu.rf_ram.memory[57][2] ;
 wire \u_cpu.rf_ram.memory[57][3] ;
 wire \u_cpu.rf_ram.memory[57][4] ;
 wire \u_cpu.rf_ram.memory[57][5] ;
 wire \u_cpu.rf_ram.memory[57][6] ;
 wire \u_cpu.rf_ram.memory[57][7] ;
 wire \u_cpu.rf_ram.memory[58][0] ;
 wire \u_cpu.rf_ram.memory[58][1] ;
 wire \u_cpu.rf_ram.memory[58][2] ;
 wire \u_cpu.rf_ram.memory[58][3] ;
 wire \u_cpu.rf_ram.memory[58][4] ;
 wire \u_cpu.rf_ram.memory[58][5] ;
 wire \u_cpu.rf_ram.memory[58][6] ;
 wire \u_cpu.rf_ram.memory[58][7] ;
 wire \u_cpu.rf_ram.memory[59][0] ;
 wire \u_cpu.rf_ram.memory[59][1] ;
 wire \u_cpu.rf_ram.memory[59][2] ;
 wire \u_cpu.rf_ram.memory[59][3] ;
 wire \u_cpu.rf_ram.memory[59][4] ;
 wire \u_cpu.rf_ram.memory[59][5] ;
 wire \u_cpu.rf_ram.memory[59][6] ;
 wire \u_cpu.rf_ram.memory[59][7] ;
 wire \u_cpu.rf_ram.memory[5][0] ;
 wire \u_cpu.rf_ram.memory[5][1] ;
 wire \u_cpu.rf_ram.memory[5][2] ;
 wire \u_cpu.rf_ram.memory[5][3] ;
 wire \u_cpu.rf_ram.memory[5][4] ;
 wire \u_cpu.rf_ram.memory[5][5] ;
 wire \u_cpu.rf_ram.memory[5][6] ;
 wire \u_cpu.rf_ram.memory[5][7] ;
 wire \u_cpu.rf_ram.memory[60][0] ;
 wire \u_cpu.rf_ram.memory[60][1] ;
 wire \u_cpu.rf_ram.memory[60][2] ;
 wire \u_cpu.rf_ram.memory[60][3] ;
 wire \u_cpu.rf_ram.memory[60][4] ;
 wire \u_cpu.rf_ram.memory[60][5] ;
 wire \u_cpu.rf_ram.memory[60][6] ;
 wire \u_cpu.rf_ram.memory[60][7] ;
 wire \u_cpu.rf_ram.memory[61][0] ;
 wire \u_cpu.rf_ram.memory[61][1] ;
 wire \u_cpu.rf_ram.memory[61][2] ;
 wire \u_cpu.rf_ram.memory[61][3] ;
 wire \u_cpu.rf_ram.memory[61][4] ;
 wire \u_cpu.rf_ram.memory[61][5] ;
 wire \u_cpu.rf_ram.memory[61][6] ;
 wire \u_cpu.rf_ram.memory[61][7] ;
 wire \u_cpu.rf_ram.memory[62][0] ;
 wire \u_cpu.rf_ram.memory[62][1] ;
 wire \u_cpu.rf_ram.memory[62][2] ;
 wire \u_cpu.rf_ram.memory[62][3] ;
 wire \u_cpu.rf_ram.memory[62][4] ;
 wire \u_cpu.rf_ram.memory[62][5] ;
 wire \u_cpu.rf_ram.memory[62][6] ;
 wire \u_cpu.rf_ram.memory[62][7] ;
 wire \u_cpu.rf_ram.memory[63][0] ;
 wire \u_cpu.rf_ram.memory[63][1] ;
 wire \u_cpu.rf_ram.memory[63][2] ;
 wire \u_cpu.rf_ram.memory[63][3] ;
 wire \u_cpu.rf_ram.memory[63][4] ;
 wire \u_cpu.rf_ram.memory[63][5] ;
 wire \u_cpu.rf_ram.memory[63][6] ;
 wire \u_cpu.rf_ram.memory[63][7] ;
 wire \u_cpu.rf_ram.memory[64][0] ;
 wire \u_cpu.rf_ram.memory[64][1] ;
 wire \u_cpu.rf_ram.memory[64][2] ;
 wire \u_cpu.rf_ram.memory[64][3] ;
 wire \u_cpu.rf_ram.memory[64][4] ;
 wire \u_cpu.rf_ram.memory[64][5] ;
 wire \u_cpu.rf_ram.memory[64][6] ;
 wire \u_cpu.rf_ram.memory[64][7] ;
 wire \u_cpu.rf_ram.memory[65][0] ;
 wire \u_cpu.rf_ram.memory[65][1] ;
 wire \u_cpu.rf_ram.memory[65][2] ;
 wire \u_cpu.rf_ram.memory[65][3] ;
 wire \u_cpu.rf_ram.memory[65][4] ;
 wire \u_cpu.rf_ram.memory[65][5] ;
 wire \u_cpu.rf_ram.memory[65][6] ;
 wire \u_cpu.rf_ram.memory[65][7] ;
 wire \u_cpu.rf_ram.memory[66][0] ;
 wire \u_cpu.rf_ram.memory[66][1] ;
 wire \u_cpu.rf_ram.memory[66][2] ;
 wire \u_cpu.rf_ram.memory[66][3] ;
 wire \u_cpu.rf_ram.memory[66][4] ;
 wire \u_cpu.rf_ram.memory[66][5] ;
 wire \u_cpu.rf_ram.memory[66][6] ;
 wire \u_cpu.rf_ram.memory[66][7] ;
 wire \u_cpu.rf_ram.memory[67][0] ;
 wire \u_cpu.rf_ram.memory[67][1] ;
 wire \u_cpu.rf_ram.memory[67][2] ;
 wire \u_cpu.rf_ram.memory[67][3] ;
 wire \u_cpu.rf_ram.memory[67][4] ;
 wire \u_cpu.rf_ram.memory[67][5] ;
 wire \u_cpu.rf_ram.memory[67][6] ;
 wire \u_cpu.rf_ram.memory[67][7] ;
 wire \u_cpu.rf_ram.memory[68][0] ;
 wire \u_cpu.rf_ram.memory[68][1] ;
 wire \u_cpu.rf_ram.memory[68][2] ;
 wire \u_cpu.rf_ram.memory[68][3] ;
 wire \u_cpu.rf_ram.memory[68][4] ;
 wire \u_cpu.rf_ram.memory[68][5] ;
 wire \u_cpu.rf_ram.memory[68][6] ;
 wire \u_cpu.rf_ram.memory[68][7] ;
 wire \u_cpu.rf_ram.memory[69][0] ;
 wire \u_cpu.rf_ram.memory[69][1] ;
 wire \u_cpu.rf_ram.memory[69][2] ;
 wire \u_cpu.rf_ram.memory[69][3] ;
 wire \u_cpu.rf_ram.memory[69][4] ;
 wire \u_cpu.rf_ram.memory[69][5] ;
 wire \u_cpu.rf_ram.memory[69][6] ;
 wire \u_cpu.rf_ram.memory[69][7] ;
 wire \u_cpu.rf_ram.memory[6][0] ;
 wire \u_cpu.rf_ram.memory[6][1] ;
 wire \u_cpu.rf_ram.memory[6][2] ;
 wire \u_cpu.rf_ram.memory[6][3] ;
 wire \u_cpu.rf_ram.memory[6][4] ;
 wire \u_cpu.rf_ram.memory[6][5] ;
 wire \u_cpu.rf_ram.memory[6][6] ;
 wire \u_cpu.rf_ram.memory[6][7] ;
 wire \u_cpu.rf_ram.memory[70][0] ;
 wire \u_cpu.rf_ram.memory[70][1] ;
 wire \u_cpu.rf_ram.memory[70][2] ;
 wire \u_cpu.rf_ram.memory[70][3] ;
 wire \u_cpu.rf_ram.memory[70][4] ;
 wire \u_cpu.rf_ram.memory[70][5] ;
 wire \u_cpu.rf_ram.memory[70][6] ;
 wire \u_cpu.rf_ram.memory[70][7] ;
 wire \u_cpu.rf_ram.memory[71][0] ;
 wire \u_cpu.rf_ram.memory[71][1] ;
 wire \u_cpu.rf_ram.memory[71][2] ;
 wire \u_cpu.rf_ram.memory[71][3] ;
 wire \u_cpu.rf_ram.memory[71][4] ;
 wire \u_cpu.rf_ram.memory[71][5] ;
 wire \u_cpu.rf_ram.memory[71][6] ;
 wire \u_cpu.rf_ram.memory[71][7] ;
 wire \u_cpu.rf_ram.memory[72][0] ;
 wire \u_cpu.rf_ram.memory[72][1] ;
 wire \u_cpu.rf_ram.memory[72][2] ;
 wire \u_cpu.rf_ram.memory[72][3] ;
 wire \u_cpu.rf_ram.memory[72][4] ;
 wire \u_cpu.rf_ram.memory[72][5] ;
 wire \u_cpu.rf_ram.memory[72][6] ;
 wire \u_cpu.rf_ram.memory[72][7] ;
 wire \u_cpu.rf_ram.memory[73][0] ;
 wire \u_cpu.rf_ram.memory[73][1] ;
 wire \u_cpu.rf_ram.memory[73][2] ;
 wire \u_cpu.rf_ram.memory[73][3] ;
 wire \u_cpu.rf_ram.memory[73][4] ;
 wire \u_cpu.rf_ram.memory[73][5] ;
 wire \u_cpu.rf_ram.memory[73][6] ;
 wire \u_cpu.rf_ram.memory[73][7] ;
 wire \u_cpu.rf_ram.memory[74][0] ;
 wire \u_cpu.rf_ram.memory[74][1] ;
 wire \u_cpu.rf_ram.memory[74][2] ;
 wire \u_cpu.rf_ram.memory[74][3] ;
 wire \u_cpu.rf_ram.memory[74][4] ;
 wire \u_cpu.rf_ram.memory[74][5] ;
 wire \u_cpu.rf_ram.memory[74][6] ;
 wire \u_cpu.rf_ram.memory[74][7] ;
 wire \u_cpu.rf_ram.memory[75][0] ;
 wire \u_cpu.rf_ram.memory[75][1] ;
 wire \u_cpu.rf_ram.memory[75][2] ;
 wire \u_cpu.rf_ram.memory[75][3] ;
 wire \u_cpu.rf_ram.memory[75][4] ;
 wire \u_cpu.rf_ram.memory[75][5] ;
 wire \u_cpu.rf_ram.memory[75][6] ;
 wire \u_cpu.rf_ram.memory[75][7] ;
 wire \u_cpu.rf_ram.memory[76][0] ;
 wire \u_cpu.rf_ram.memory[76][1] ;
 wire \u_cpu.rf_ram.memory[76][2] ;
 wire \u_cpu.rf_ram.memory[76][3] ;
 wire \u_cpu.rf_ram.memory[76][4] ;
 wire \u_cpu.rf_ram.memory[76][5] ;
 wire \u_cpu.rf_ram.memory[76][6] ;
 wire \u_cpu.rf_ram.memory[76][7] ;
 wire \u_cpu.rf_ram.memory[77][0] ;
 wire \u_cpu.rf_ram.memory[77][1] ;
 wire \u_cpu.rf_ram.memory[77][2] ;
 wire \u_cpu.rf_ram.memory[77][3] ;
 wire \u_cpu.rf_ram.memory[77][4] ;
 wire \u_cpu.rf_ram.memory[77][5] ;
 wire \u_cpu.rf_ram.memory[77][6] ;
 wire \u_cpu.rf_ram.memory[77][7] ;
 wire \u_cpu.rf_ram.memory[78][0] ;
 wire \u_cpu.rf_ram.memory[78][1] ;
 wire \u_cpu.rf_ram.memory[78][2] ;
 wire \u_cpu.rf_ram.memory[78][3] ;
 wire \u_cpu.rf_ram.memory[78][4] ;
 wire \u_cpu.rf_ram.memory[78][5] ;
 wire \u_cpu.rf_ram.memory[78][6] ;
 wire \u_cpu.rf_ram.memory[78][7] ;
 wire \u_cpu.rf_ram.memory[79][0] ;
 wire \u_cpu.rf_ram.memory[79][1] ;
 wire \u_cpu.rf_ram.memory[79][2] ;
 wire \u_cpu.rf_ram.memory[79][3] ;
 wire \u_cpu.rf_ram.memory[79][4] ;
 wire \u_cpu.rf_ram.memory[79][5] ;
 wire \u_cpu.rf_ram.memory[79][6] ;
 wire \u_cpu.rf_ram.memory[79][7] ;
 wire \u_cpu.rf_ram.memory[7][0] ;
 wire \u_cpu.rf_ram.memory[7][1] ;
 wire \u_cpu.rf_ram.memory[7][2] ;
 wire \u_cpu.rf_ram.memory[7][3] ;
 wire \u_cpu.rf_ram.memory[7][4] ;
 wire \u_cpu.rf_ram.memory[7][5] ;
 wire \u_cpu.rf_ram.memory[7][6] ;
 wire \u_cpu.rf_ram.memory[7][7] ;
 wire \u_cpu.rf_ram.memory[80][0] ;
 wire \u_cpu.rf_ram.memory[80][1] ;
 wire \u_cpu.rf_ram.memory[80][2] ;
 wire \u_cpu.rf_ram.memory[80][3] ;
 wire \u_cpu.rf_ram.memory[80][4] ;
 wire \u_cpu.rf_ram.memory[80][5] ;
 wire \u_cpu.rf_ram.memory[80][6] ;
 wire \u_cpu.rf_ram.memory[80][7] ;
 wire \u_cpu.rf_ram.memory[81][0] ;
 wire \u_cpu.rf_ram.memory[81][1] ;
 wire \u_cpu.rf_ram.memory[81][2] ;
 wire \u_cpu.rf_ram.memory[81][3] ;
 wire \u_cpu.rf_ram.memory[81][4] ;
 wire \u_cpu.rf_ram.memory[81][5] ;
 wire \u_cpu.rf_ram.memory[81][6] ;
 wire \u_cpu.rf_ram.memory[81][7] ;
 wire \u_cpu.rf_ram.memory[82][0] ;
 wire \u_cpu.rf_ram.memory[82][1] ;
 wire \u_cpu.rf_ram.memory[82][2] ;
 wire \u_cpu.rf_ram.memory[82][3] ;
 wire \u_cpu.rf_ram.memory[82][4] ;
 wire \u_cpu.rf_ram.memory[82][5] ;
 wire \u_cpu.rf_ram.memory[82][6] ;
 wire \u_cpu.rf_ram.memory[82][7] ;
 wire \u_cpu.rf_ram.memory[83][0] ;
 wire \u_cpu.rf_ram.memory[83][1] ;
 wire \u_cpu.rf_ram.memory[83][2] ;
 wire \u_cpu.rf_ram.memory[83][3] ;
 wire \u_cpu.rf_ram.memory[83][4] ;
 wire \u_cpu.rf_ram.memory[83][5] ;
 wire \u_cpu.rf_ram.memory[83][6] ;
 wire \u_cpu.rf_ram.memory[83][7] ;
 wire \u_cpu.rf_ram.memory[84][0] ;
 wire \u_cpu.rf_ram.memory[84][1] ;
 wire \u_cpu.rf_ram.memory[84][2] ;
 wire \u_cpu.rf_ram.memory[84][3] ;
 wire \u_cpu.rf_ram.memory[84][4] ;
 wire \u_cpu.rf_ram.memory[84][5] ;
 wire \u_cpu.rf_ram.memory[84][6] ;
 wire \u_cpu.rf_ram.memory[84][7] ;
 wire \u_cpu.rf_ram.memory[85][0] ;
 wire \u_cpu.rf_ram.memory[85][1] ;
 wire \u_cpu.rf_ram.memory[85][2] ;
 wire \u_cpu.rf_ram.memory[85][3] ;
 wire \u_cpu.rf_ram.memory[85][4] ;
 wire \u_cpu.rf_ram.memory[85][5] ;
 wire \u_cpu.rf_ram.memory[85][6] ;
 wire \u_cpu.rf_ram.memory[85][7] ;
 wire \u_cpu.rf_ram.memory[86][0] ;
 wire \u_cpu.rf_ram.memory[86][1] ;
 wire \u_cpu.rf_ram.memory[86][2] ;
 wire \u_cpu.rf_ram.memory[86][3] ;
 wire \u_cpu.rf_ram.memory[86][4] ;
 wire \u_cpu.rf_ram.memory[86][5] ;
 wire \u_cpu.rf_ram.memory[86][6] ;
 wire \u_cpu.rf_ram.memory[86][7] ;
 wire \u_cpu.rf_ram.memory[87][0] ;
 wire \u_cpu.rf_ram.memory[87][1] ;
 wire \u_cpu.rf_ram.memory[87][2] ;
 wire \u_cpu.rf_ram.memory[87][3] ;
 wire \u_cpu.rf_ram.memory[87][4] ;
 wire \u_cpu.rf_ram.memory[87][5] ;
 wire \u_cpu.rf_ram.memory[87][6] ;
 wire \u_cpu.rf_ram.memory[87][7] ;
 wire \u_cpu.rf_ram.memory[88][0] ;
 wire \u_cpu.rf_ram.memory[88][1] ;
 wire \u_cpu.rf_ram.memory[88][2] ;
 wire \u_cpu.rf_ram.memory[88][3] ;
 wire \u_cpu.rf_ram.memory[88][4] ;
 wire \u_cpu.rf_ram.memory[88][5] ;
 wire \u_cpu.rf_ram.memory[88][6] ;
 wire \u_cpu.rf_ram.memory[88][7] ;
 wire \u_cpu.rf_ram.memory[89][0] ;
 wire \u_cpu.rf_ram.memory[89][1] ;
 wire \u_cpu.rf_ram.memory[89][2] ;
 wire \u_cpu.rf_ram.memory[89][3] ;
 wire \u_cpu.rf_ram.memory[89][4] ;
 wire \u_cpu.rf_ram.memory[89][5] ;
 wire \u_cpu.rf_ram.memory[89][6] ;
 wire \u_cpu.rf_ram.memory[89][7] ;
 wire \u_cpu.rf_ram.memory[8][0] ;
 wire \u_cpu.rf_ram.memory[8][1] ;
 wire \u_cpu.rf_ram.memory[8][2] ;
 wire \u_cpu.rf_ram.memory[8][3] ;
 wire \u_cpu.rf_ram.memory[8][4] ;
 wire \u_cpu.rf_ram.memory[8][5] ;
 wire \u_cpu.rf_ram.memory[8][6] ;
 wire \u_cpu.rf_ram.memory[8][7] ;
 wire \u_cpu.rf_ram.memory[90][0] ;
 wire \u_cpu.rf_ram.memory[90][1] ;
 wire \u_cpu.rf_ram.memory[90][2] ;
 wire \u_cpu.rf_ram.memory[90][3] ;
 wire \u_cpu.rf_ram.memory[90][4] ;
 wire \u_cpu.rf_ram.memory[90][5] ;
 wire \u_cpu.rf_ram.memory[90][6] ;
 wire \u_cpu.rf_ram.memory[90][7] ;
 wire \u_cpu.rf_ram.memory[91][0] ;
 wire \u_cpu.rf_ram.memory[91][1] ;
 wire \u_cpu.rf_ram.memory[91][2] ;
 wire \u_cpu.rf_ram.memory[91][3] ;
 wire \u_cpu.rf_ram.memory[91][4] ;
 wire \u_cpu.rf_ram.memory[91][5] ;
 wire \u_cpu.rf_ram.memory[91][6] ;
 wire \u_cpu.rf_ram.memory[91][7] ;
 wire \u_cpu.rf_ram.memory[92][0] ;
 wire \u_cpu.rf_ram.memory[92][1] ;
 wire \u_cpu.rf_ram.memory[92][2] ;
 wire \u_cpu.rf_ram.memory[92][3] ;
 wire \u_cpu.rf_ram.memory[92][4] ;
 wire \u_cpu.rf_ram.memory[92][5] ;
 wire \u_cpu.rf_ram.memory[92][6] ;
 wire \u_cpu.rf_ram.memory[92][7] ;
 wire \u_cpu.rf_ram.memory[93][0] ;
 wire \u_cpu.rf_ram.memory[93][1] ;
 wire \u_cpu.rf_ram.memory[93][2] ;
 wire \u_cpu.rf_ram.memory[93][3] ;
 wire \u_cpu.rf_ram.memory[93][4] ;
 wire \u_cpu.rf_ram.memory[93][5] ;
 wire \u_cpu.rf_ram.memory[93][6] ;
 wire \u_cpu.rf_ram.memory[93][7] ;
 wire \u_cpu.rf_ram.memory[94][0] ;
 wire \u_cpu.rf_ram.memory[94][1] ;
 wire \u_cpu.rf_ram.memory[94][2] ;
 wire \u_cpu.rf_ram.memory[94][3] ;
 wire \u_cpu.rf_ram.memory[94][4] ;
 wire \u_cpu.rf_ram.memory[94][5] ;
 wire \u_cpu.rf_ram.memory[94][6] ;
 wire \u_cpu.rf_ram.memory[94][7] ;
 wire \u_cpu.rf_ram.memory[95][0] ;
 wire \u_cpu.rf_ram.memory[95][1] ;
 wire \u_cpu.rf_ram.memory[95][2] ;
 wire \u_cpu.rf_ram.memory[95][3] ;
 wire \u_cpu.rf_ram.memory[95][4] ;
 wire \u_cpu.rf_ram.memory[95][5] ;
 wire \u_cpu.rf_ram.memory[95][6] ;
 wire \u_cpu.rf_ram.memory[95][7] ;
 wire \u_cpu.rf_ram.memory[96][0] ;
 wire \u_cpu.rf_ram.memory[96][1] ;
 wire \u_cpu.rf_ram.memory[96][2] ;
 wire \u_cpu.rf_ram.memory[96][3] ;
 wire \u_cpu.rf_ram.memory[96][4] ;
 wire \u_cpu.rf_ram.memory[96][5] ;
 wire \u_cpu.rf_ram.memory[96][6] ;
 wire \u_cpu.rf_ram.memory[96][7] ;
 wire \u_cpu.rf_ram.memory[97][0] ;
 wire \u_cpu.rf_ram.memory[97][1] ;
 wire \u_cpu.rf_ram.memory[97][2] ;
 wire \u_cpu.rf_ram.memory[97][3] ;
 wire \u_cpu.rf_ram.memory[97][4] ;
 wire \u_cpu.rf_ram.memory[97][5] ;
 wire \u_cpu.rf_ram.memory[97][6] ;
 wire \u_cpu.rf_ram.memory[97][7] ;
 wire \u_cpu.rf_ram.memory[98][0] ;
 wire \u_cpu.rf_ram.memory[98][1] ;
 wire \u_cpu.rf_ram.memory[98][2] ;
 wire \u_cpu.rf_ram.memory[98][3] ;
 wire \u_cpu.rf_ram.memory[98][4] ;
 wire \u_cpu.rf_ram.memory[98][5] ;
 wire \u_cpu.rf_ram.memory[98][6] ;
 wire \u_cpu.rf_ram.memory[98][7] ;
 wire \u_cpu.rf_ram.memory[99][0] ;
 wire \u_cpu.rf_ram.memory[99][1] ;
 wire \u_cpu.rf_ram.memory[99][2] ;
 wire \u_cpu.rf_ram.memory[99][3] ;
 wire \u_cpu.rf_ram.memory[99][4] ;
 wire \u_cpu.rf_ram.memory[99][5] ;
 wire \u_cpu.rf_ram.memory[99][6] ;
 wire \u_cpu.rf_ram.memory[99][7] ;
 wire \u_cpu.rf_ram.memory[9][0] ;
 wire \u_cpu.rf_ram.memory[9][1] ;
 wire \u_cpu.rf_ram.memory[9][2] ;
 wire \u_cpu.rf_ram.memory[9][3] ;
 wire \u_cpu.rf_ram.memory[9][4] ;
 wire \u_cpu.rf_ram.memory[9][5] ;
 wire \u_cpu.rf_ram.memory[9][6] ;
 wire \u_cpu.rf_ram.memory[9][7] ;
 wire \u_cpu.rf_ram.rdata[0] ;
 wire \u_cpu.rf_ram.rdata[1] ;
 wire \u_cpu.rf_ram.rdata[2] ;
 wire \u_cpu.rf_ram.rdata[3] ;
 wire \u_cpu.rf_ram.rdata[4] ;
 wire \u_cpu.rf_ram.rdata[5] ;
 wire \u_cpu.rf_ram.rdata[6] ;
 wire \u_cpu.rf_ram.rdata[7] ;
 wire \u_cpu.rf_ram.regzero ;
 wire \u_cpu.rf_ram_if.genblk1.wtrig0_r ;
 wire \u_cpu.rf_ram_if.rcnt[0] ;
 wire \u_cpu.rf_ram_if.rcnt[1] ;
 wire \u_cpu.rf_ram_if.rcnt[2] ;
 wire \u_cpu.rf_ram_if.rdata0[1] ;
 wire \u_cpu.rf_ram_if.rdata0[2] ;
 wire \u_cpu.rf_ram_if.rdata0[3] ;
 wire \u_cpu.rf_ram_if.rdata0[4] ;
 wire \u_cpu.rf_ram_if.rdata0[5] ;
 wire \u_cpu.rf_ram_if.rdata0[6] ;
 wire \u_cpu.rf_ram_if.rdata0[7] ;
 wire \u_cpu.rf_ram_if.rdata1[0] ;
 wire \u_cpu.rf_ram_if.rdata1[1] ;
 wire \u_cpu.rf_ram_if.rdata1[2] ;
 wire \u_cpu.rf_ram_if.rdata1[3] ;
 wire \u_cpu.rf_ram_if.rdata1[4] ;
 wire \u_cpu.rf_ram_if.rdata1[5] ;
 wire \u_cpu.rf_ram_if.rdata1[6] ;
 wire \u_cpu.rf_ram_if.rgnt ;
 wire \u_cpu.rf_ram_if.rreq_r ;
 wire \u_cpu.rf_ram_if.rtrig0 ;
 wire \u_cpu.rf_ram_if.rtrig1 ;
 wire \u_cpu.rf_ram_if.wdata0_r[0] ;
 wire \u_cpu.rf_ram_if.wdata0_r[1] ;
 wire \u_cpu.rf_ram_if.wdata0_r[2] ;
 wire \u_cpu.rf_ram_if.wdata0_r[3] ;
 wire \u_cpu.rf_ram_if.wdata0_r[4] ;
 wire \u_cpu.rf_ram_if.wdata0_r[5] ;
 wire \u_cpu.rf_ram_if.wdata0_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \u_cpu.rf_ram_if.wdata1_r[2] ;
 wire \u_cpu.rf_ram_if.wdata1_r[3] ;
 wire \u_cpu.rf_ram_if.wdata1_r[4] ;
 wire \u_cpu.rf_ram_if.wdata1_r[5] ;
 wire \u_cpu.rf_ram_if.wdata1_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[7] ;
 wire \u_cpu.rf_ram_if.wen0_r ;
 wire \u_cpu.rf_ram_if.wen1_r ;
 wire \u_cpu.rf_ram_if.wtrig0 ;
 wire \u_scanchain_local.data_out ;
 wire \u_scanchain_local.module_data_in[34] ;
 wire \u_scanchain_local.module_data_in[35] ;
 wire \u_scanchain_local.module_data_in[36] ;
 wire \u_scanchain_local.module_data_in[37] ;
 wire \u_scanchain_local.module_data_in[38] ;
 wire \u_scanchain_local.module_data_in[39] ;
 wire \u_scanchain_local.module_data_in[40] ;
 wire \u_scanchain_local.module_data_in[41] ;
 wire \u_scanchain_local.module_data_in[42] ;
 wire \u_scanchain_local.module_data_in[43] ;
 wire \u_scanchain_local.module_data_in[44] ;
 wire \u_scanchain_local.module_data_in[45] ;
 wire \u_scanchain_local.module_data_in[46] ;
 wire \u_scanchain_local.module_data_in[47] ;
 wire \u_scanchain_local.module_data_in[48] ;
 wire \u_scanchain_local.module_data_in[49] ;
 wire \u_scanchain_local.module_data_in[50] ;
 wire \u_scanchain_local.module_data_in[51] ;
 wire \u_scanchain_local.module_data_in[52] ;
 wire \u_scanchain_local.module_data_in[53] ;
 wire \u_scanchain_local.module_data_in[54] ;
 wire \u_scanchain_local.module_data_in[55] ;
 wire \u_scanchain_local.module_data_in[56] ;
 wire \u_scanchain_local.module_data_in[57] ;
 wire \u_scanchain_local.module_data_in[58] ;
 wire \u_scanchain_local.module_data_in[59] ;
 wire \u_scanchain_local.module_data_in[60] ;
 wire \u_scanchain_local.module_data_in[61] ;
 wire \u_scanchain_local.module_data_in[62] ;
 wire \u_scanchain_local.module_data_in[63] ;
 wire \u_scanchain_local.module_data_in[64] ;
 wire \u_scanchain_local.module_data_in[65] ;
 wire \u_scanchain_local.module_data_in[66] ;
 wire \u_scanchain_local.module_data_in[67] ;
 wire \u_scanchain_local.module_data_in[68] ;
 wire \u_scanchain_local.module_data_in[69] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05784_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05785_ (.A1(_01436_),
    .A2(\u_cpu.rf_ram_if.rcnt[2] ),
    .A3(\u_cpu.rf_ram_if.rcnt[1] ),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05786_ (.I(_01437_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05787_ (.I(_01438_),
    .Z(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05788_ (.I(\u_cpu.cpu.csr_imm ),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05789_ (.I(_01437_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05790_ (.I(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05791_ (.A1(\u_cpu.cpu.decode.co_mem_word ),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .A3(\u_cpu.cpu.csr_d_sel ),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05792_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05793_ (.I(\u_cpu.cpu.branch_op ),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05794_ (.A1(_01443_),
    .A2(_01444_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05795_ (.A1(_01442_),
    .A2(_01445_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05796_ (.I(_01446_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05797_ (.I(\u_cpu.cpu.decode.op21 ),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05798_ (.I(\u_cpu.cpu.decode.co_ebreak ),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05799_ (.A1(_01448_),
    .A2(\u_cpu.cpu.decode.op26 ),
    .B(_01449_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05800_ (.I(\u_cpu.cpu.decode.co_mem_word ),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05801_ (.I(\u_cpu.cpu.csr_d_sel ),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05802_ (.A1(_01451_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .A3(_01452_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05803_ (.A1(_01453_),
    .A2(_01445_),
    .B(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .C(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05804_ (.A1(_01447_),
    .A2(_01450_),
    .B(_01454_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05805_ (.A1(_01441_),
    .A2(_01455_),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05806_ (.I(\u_cpu.cpu.decode.op26 ),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05807_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05808_ (.A1(_01447_),
    .A2(_01450_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05809_ (.A1(_01443_),
    .A2(_01444_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05810_ (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05811_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01442_),
    .A3(_01460_),
    .B(_01461_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05812_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_01462_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05813_ (.A1(_01458_),
    .A2(_01459_),
    .B(_01438_),
    .C(_01463_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05814_ (.A1(_01456_),
    .A2(_01464_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05815_ (.A1(_01439_),
    .A2(_01440_),
    .B(_01465_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05816_ (.I(_01466_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05817_ (.I(_01467_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05818_ (.I(_01468_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05819_ (.A1(\u_cpu.rf_ram_if.rtrig0 ),
    .A2(_01455_),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05820_ (.I(_01440_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05821_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_01471_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05822_ (.A1(_01440_),
    .A2(_01455_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05823_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_01473_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05824_ (.A1(_01472_),
    .A2(_01474_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05825_ (.A1(_01470_),
    .A2(_01475_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05826_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05827_ (.I(\u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05828_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_01449_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05829_ (.A1(_01448_),
    .A2(_01442_),
    .A3(_01460_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05830_ (.A1(_01440_),
    .A2(_01480_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _05831_ (.A1(_01478_),
    .A2(_01455_),
    .B1(_01479_),
    .B2(_01447_),
    .C(_01481_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05832_ (.A1(_01477_),
    .A2(_01482_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05833_ (.I(_01483_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05834_ (.I(_01484_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05835_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_01440_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05836_ (.A1(\u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_01473_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05837_ (.A1(_01486_),
    .A2(_01487_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05838_ (.I(_01488_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05839_ (.I(_01489_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05840_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_01471_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05841_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_01473_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05842_ (.A1(_01491_),
    .A2(_01492_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05843_ (.I(_01493_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05844_ (.A1(_01476_),
    .A2(_01485_),
    .A3(_01490_),
    .A4(_01494_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05845_ (.A1(_01469_),
    .A2(_01495_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05846_ (.I(_01471_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05847_ (.I(_01496_),
    .ZN(\u_cpu.rf_ram_if.wtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05848_ (.I(_01476_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05849_ (.A1(_01491_),
    .A2(_01492_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05850_ (.I(_01498_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05851_ (.I(_01467_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05852_ (.I(\u_cpu.raddr[0] ),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05853_ (.I(_01501_),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05854_ (.I(_01502_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05855_ (.I(_01503_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05856_ (.I(\u_cpu.raddr[1] ),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05857_ (.I(_01505_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05858_ (.I(_01506_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05859_ (.I0(\u_cpu.rf_ram.memory[28][0] ),
    .I1(\u_cpu.rf_ram.memory[29][0] ),
    .I2(\u_cpu.rf_ram.memory[30][0] ),
    .I3(\u_cpu.rf_ram.memory[31][0] ),
    .S0(_01504_),
    .S1(_01507_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05860_ (.A1(_01500_),
    .A2(_01508_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05861_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(\u_cpu.rf_ram_if.rtrig0 ),
    .B1(_01456_),
    .B2(_01464_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05862_ (.I(_01510_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05863_ (.I(_01511_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05864_ (.I(_01512_),
    .Z(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05865_ (.I(\u_cpu.raddr[0] ),
    .Z(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05866_ (.I(_01514_),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05867_ (.I(_01515_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05868_ (.I(_01505_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05869_ (.I(_01517_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05870_ (.I0(\u_cpu.rf_ram.memory[24][0] ),
    .I1(\u_cpu.rf_ram.memory[25][0] ),
    .I2(\u_cpu.rf_ram.memory[26][0] ),
    .I3(\u_cpu.rf_ram.memory[27][0] ),
    .S0(_01516_),
    .S1(_01518_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05871_ (.I(_01483_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05872_ (.I(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05873_ (.A1(_01513_),
    .A2(_01519_),
    .B(_01521_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05874_ (.I(_01467_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05875_ (.I(_01503_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05876_ (.I(_01506_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05877_ (.I0(\u_cpu.rf_ram.memory[20][0] ),
    .I1(\u_cpu.rf_ram.memory[21][0] ),
    .I2(\u_cpu.rf_ram.memory[22][0] ),
    .I3(\u_cpu.rf_ram.memory[23][0] ),
    .S0(_01524_),
    .S1(_01525_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05878_ (.A1(_01523_),
    .A2(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05879_ (.I(_01512_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05880_ (.I(_01515_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05881_ (.I(_01517_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05882_ (.I0(\u_cpu.rf_ram.memory[16][0] ),
    .I1(\u_cpu.rf_ram.memory[17][0] ),
    .I2(\u_cpu.rf_ram.memory[18][0] ),
    .I3(\u_cpu.rf_ram.memory[19][0] ),
    .S0(_01529_),
    .S1(_01530_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05883_ (.A1(_01477_),
    .A2(_01482_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05884_ (.I(_01532_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05885_ (.I(_01533_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05886_ (.A1(_01528_),
    .A2(_01531_),
    .B(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05887_ (.A1(_01509_),
    .A2(_01522_),
    .B1(_01527_),
    .B2(_01535_),
    .C(_01490_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05888_ (.I(_01466_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05889_ (.I(_01537_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05890_ (.I(_01538_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05891_ (.I(_01514_),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05892_ (.I(_01540_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05893_ (.I(_01541_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05894_ (.I(_01505_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05895_ (.I(_01543_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05896_ (.I0(\u_cpu.rf_ram.memory[4][0] ),
    .I1(\u_cpu.rf_ram.memory[5][0] ),
    .I2(\u_cpu.rf_ram.memory[6][0] ),
    .I3(\u_cpu.rf_ram.memory[7][0] ),
    .S0(_01542_),
    .S1(_01544_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05897_ (.A1(_01539_),
    .A2(_01545_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05898_ (.I(_01512_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05899_ (.I(_01501_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05900_ (.I(_01548_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05901_ (.I(_01549_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05902_ (.I(\u_cpu.raddr[1] ),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05903_ (.I(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05904_ (.I(_01552_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05905_ (.I0(\u_cpu.rf_ram.memory[0][0] ),
    .I1(\u_cpu.rf_ram.memory[1][0] ),
    .I2(\u_cpu.rf_ram.memory[2][0] ),
    .I3(\u_cpu.rf_ram.memory[3][0] ),
    .S0(_01550_),
    .S1(_01553_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05906_ (.I(_01532_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05907_ (.I(_01555_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05908_ (.A1(_01547_),
    .A2(_01554_),
    .B(_01556_),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05909_ (.I(_01510_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05910_ (.I(_01558_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05911_ (.I(_01559_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05912_ (.I(_01503_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05913_ (.I(_01551_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05914_ (.I(_01562_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05915_ (.I(_01563_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05916_ (.I0(\u_cpu.rf_ram.memory[8][0] ),
    .I1(\u_cpu.rf_ram.memory[9][0] ),
    .I2(\u_cpu.rf_ram.memory[10][0] ),
    .I3(\u_cpu.rf_ram.memory[11][0] ),
    .S0(_01561_),
    .S1(_01564_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05917_ (.A1(_01560_),
    .A2(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05918_ (.I(_01467_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05919_ (.I(_01501_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05920_ (.I(_01568_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05921_ (.I(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05922_ (.I(_01505_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05923_ (.I(_01571_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05924_ (.I0(\u_cpu.rf_ram.memory[12][0] ),
    .I1(\u_cpu.rf_ram.memory[13][0] ),
    .I2(\u_cpu.rf_ram.memory[14][0] ),
    .I3(\u_cpu.rf_ram.memory[15][0] ),
    .S0(_01570_),
    .S1(_01572_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05925_ (.I(_01484_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05926_ (.A1(_01567_),
    .A2(_01573_),
    .B(_01574_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05927_ (.A1(_01486_),
    .A2(_01487_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05928_ (.I(_01576_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05929_ (.I(_01577_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05930_ (.A1(_01546_),
    .A2(_01557_),
    .B1(_01566_),
    .B2(_01575_),
    .C(_01578_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05931_ (.I(_01493_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05932_ (.I(_01466_),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05933_ (.I(_01581_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05934_ (.I(_01514_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05935_ (.I(_01583_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05936_ (.I(_01551_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05937_ (.I(_01585_),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05938_ (.I0(\u_cpu.rf_ram.memory[36][0] ),
    .I1(\u_cpu.rf_ram.memory[37][0] ),
    .I2(\u_cpu.rf_ram.memory[38][0] ),
    .I3(\u_cpu.rf_ram.memory[39][0] ),
    .S0(_01584_),
    .S1(_01586_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05939_ (.A1(_01582_),
    .A2(_01587_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05940_ (.I(_01511_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05941_ (.I(_01548_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05942_ (.I(\u_cpu.raddr[1] ),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05943_ (.I(_01591_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05944_ (.I(_01592_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05945_ (.I0(\u_cpu.rf_ram.memory[32][0] ),
    .I1(\u_cpu.rf_ram.memory[33][0] ),
    .I2(\u_cpu.rf_ram.memory[34][0] ),
    .I3(\u_cpu.rf_ram.memory[35][0] ),
    .S0(_01590_),
    .S1(_01593_),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05946_ (.I(_01532_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05947_ (.I(_01595_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05948_ (.A1(_01589_),
    .A2(_01594_),
    .B(_01596_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05949_ (.I(_01510_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05950_ (.I(_01598_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05951_ (.I(_01551_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05952_ (.I(_01600_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05953_ (.I0(\u_cpu.rf_ram.memory[40][0] ),
    .I1(\u_cpu.rf_ram.memory[41][0] ),
    .I2(\u_cpu.rf_ram.memory[42][0] ),
    .I3(\u_cpu.rf_ram.memory[43][0] ),
    .S0(_01569_),
    .S1(_01601_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05954_ (.A1(_01599_),
    .A2(_01602_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05955_ (.I(_01537_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05956_ (.I(_01501_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05957_ (.I(_01605_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05958_ (.I(_01591_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05959_ (.I(_01607_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05960_ (.I0(\u_cpu.rf_ram.memory[44][0] ),
    .I1(\u_cpu.rf_ram.memory[45][0] ),
    .I2(\u_cpu.rf_ram.memory[46][0] ),
    .I3(\u_cpu.rf_ram.memory[47][0] ),
    .S0(_01606_),
    .S1(_01608_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05961_ (.I(_01483_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05962_ (.I(_01610_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05963_ (.A1(_01604_),
    .A2(_01609_),
    .B(_01611_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05964_ (.I(_01576_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05965_ (.A1(_01588_),
    .A2(_01597_),
    .B1(_01603_),
    .B2(_01612_),
    .C(_01613_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05966_ (.I(_01581_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05967_ (.I(_01514_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05968_ (.I(_01616_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05969_ (.I(_01551_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05970_ (.I(_01618_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05971_ (.I0(\u_cpu.rf_ram.memory[60][0] ),
    .I1(\u_cpu.rf_ram.memory[61][0] ),
    .I2(\u_cpu.rf_ram.memory[62][0] ),
    .I3(\u_cpu.rf_ram.memory[63][0] ),
    .S0(_01617_),
    .S1(_01619_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05972_ (.A1(_01615_),
    .A2(_01620_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05973_ (.I(_01511_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05974_ (.I(_01548_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05975_ (.I(_01592_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05976_ (.I0(\u_cpu.rf_ram.memory[56][0] ),
    .I1(\u_cpu.rf_ram.memory[57][0] ),
    .I2(\u_cpu.rf_ram.memory[58][0] ),
    .I3(\u_cpu.rf_ram.memory[59][0] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05977_ (.I(_01483_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05978_ (.A1(_01622_),
    .A2(_01625_),
    .B(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05979_ (.I(_01466_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05980_ (.I(_01628_),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05981_ (.I(_01583_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05982_ (.I(_01600_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05983_ (.I0(\u_cpu.rf_ram.memory[52][0] ),
    .I1(\u_cpu.rf_ram.memory[53][0] ),
    .I2(\u_cpu.rf_ram.memory[54][0] ),
    .I3(\u_cpu.rf_ram.memory[55][0] ),
    .S0(_01630_),
    .S1(_01631_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05984_ (.A1(_01629_),
    .A2(_01632_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05985_ (.I(_01598_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05986_ (.I(_01501_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05987_ (.I(_01635_),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05988_ (.I(_01591_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05989_ (.I(_01637_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05990_ (.I0(\u_cpu.rf_ram.memory[48][0] ),
    .I1(\u_cpu.rf_ram.memory[49][0] ),
    .I2(\u_cpu.rf_ram.memory[50][0] ),
    .I3(\u_cpu.rf_ram.memory[51][0] ),
    .S0(_01636_),
    .S1(_01638_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05991_ (.I(_01595_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05992_ (.A1(_01634_),
    .A2(_01639_),
    .B(_01640_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05993_ (.I(_01488_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05994_ (.A1(_01621_),
    .A2(_01627_),
    .B1(_01633_),
    .B2(_01641_),
    .C(_01642_),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05995_ (.A1(_01580_),
    .A2(_01614_),
    .A3(_01643_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05996_ (.A1(_01499_),
    .A2(_01536_),
    .A3(_01579_),
    .B(_01644_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05997_ (.I(_01628_),
    .Z(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05998_ (.I(_01568_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05999_ (.I(_01600_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06000_ (.I0(\u_cpu.rf_ram.memory[100][0] ),
    .I1(\u_cpu.rf_ram.memory[101][0] ),
    .I2(\u_cpu.rf_ram.memory[102][0] ),
    .I3(\u_cpu.rf_ram.memory[103][0] ),
    .S0(_01647_),
    .S1(_01648_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06001_ (.A1(_01646_),
    .A2(_01649_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06002_ (.I(_01511_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06003_ (.I(_01548_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06004_ (.I0(\u_cpu.rf_ram.memory[96][0] ),
    .I1(\u_cpu.rf_ram.memory[97][0] ),
    .I2(\u_cpu.rf_ram.memory[98][0] ),
    .I3(\u_cpu.rf_ram.memory[99][0] ),
    .S0(_01652_),
    .S1(_01552_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06005_ (.I(_01595_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06006_ (.A1(_01651_),
    .A2(_01653_),
    .B(_01654_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06007_ (.I(_01628_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06008_ (.I0(\u_cpu.rf_ram.memory[108][0] ),
    .I1(\u_cpu.rf_ram.memory[109][0] ),
    .I2(\u_cpu.rf_ram.memory[110][0] ),
    .I3(\u_cpu.rf_ram.memory[111][0] ),
    .S0(_01549_),
    .S1(_01563_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06009_ (.A1(_01656_),
    .A2(_01657_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06010_ (.I(_01510_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06011_ (.I(_01659_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06012_ (.I(_01605_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06013_ (.I0(\u_cpu.rf_ram.memory[104][0] ),
    .I1(\u_cpu.rf_ram.memory[105][0] ),
    .I2(\u_cpu.rf_ram.memory[106][0] ),
    .I3(\u_cpu.rf_ram.memory[107][0] ),
    .S0(_01661_),
    .S1(_01571_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06014_ (.I(_01610_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06015_ (.A1(_01660_),
    .A2(_01662_),
    .B(_01663_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06016_ (.I(_01576_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06017_ (.A1(_01650_),
    .A2(_01655_),
    .B1(_01658_),
    .B2(_01664_),
    .C(_01665_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06018_ (.I(_01581_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06019_ (.I(_01616_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06020_ (.I(_01618_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06021_ (.I0(\u_cpu.rf_ram.memory[124][0] ),
    .I1(\u_cpu.rf_ram.memory[125][0] ),
    .I2(\u_cpu.rf_ram.memory[126][0] ),
    .I3(\u_cpu.rf_ram.memory[127][0] ),
    .S0(_01668_),
    .S1(_01669_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06022_ (.A1(_01667_),
    .A2(_01670_),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06023_ (.I(_01659_),
    .Z(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06024_ (.I(_01605_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06025_ (.I(_01607_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06026_ (.I0(\u_cpu.rf_ram.memory[120][0] ),
    .I1(\u_cpu.rf_ram.memory[121][0] ),
    .I2(\u_cpu.rf_ram.memory[122][0] ),
    .I3(\u_cpu.rf_ram.memory[123][0] ),
    .S0(_01673_),
    .S1(_01674_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06027_ (.I(_01610_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06028_ (.A1(_01672_),
    .A2(_01675_),
    .B(_01676_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06029_ (.I(_01598_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06030_ (.I(_01583_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06031_ (.I(_01585_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06032_ (.I0(\u_cpu.rf_ram.memory[112][0] ),
    .I1(\u_cpu.rf_ram.memory[113][0] ),
    .I2(\u_cpu.rf_ram.memory[114][0] ),
    .I3(\u_cpu.rf_ram.memory[115][0] ),
    .S0(_01679_),
    .S1(_01680_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06033_ (.A1(_01678_),
    .A2(_01681_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06034_ (.I(_01537_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06035_ (.I(_01635_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06036_ (.I(_01637_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06037_ (.I0(\u_cpu.rf_ram.memory[116][0] ),
    .I1(\u_cpu.rf_ram.memory[117][0] ),
    .I2(\u_cpu.rf_ram.memory[118][0] ),
    .I3(\u_cpu.rf_ram.memory[119][0] ),
    .S0(_01684_),
    .S1(_01685_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06038_ (.I(_01595_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06039_ (.A1(_01683_),
    .A2(_01686_),
    .B(_01687_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06040_ (.I(_01488_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06041_ (.A1(_01671_),
    .A2(_01677_),
    .B1(_01682_),
    .B2(_01688_),
    .C(_01689_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06042_ (.A1(_01494_),
    .A2(_01666_),
    .A3(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06043_ (.I(_01498_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06044_ (.I(_01581_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06045_ (.I(_01540_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06046_ (.I(_01618_),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06047_ (.I0(\u_cpu.rf_ram.memory[92][0] ),
    .I1(\u_cpu.rf_ram.memory[93][0] ),
    .I2(\u_cpu.rf_ram.memory[94][0] ),
    .I3(\u_cpu.rf_ram.memory[95][0] ),
    .S0(_01694_),
    .S1(_01695_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06048_ (.A1(_01693_),
    .A2(_01696_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06049_ (.I(_01659_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06050_ (.I(_01635_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06051_ (.I(_01607_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06052_ (.I0(\u_cpu.rf_ram.memory[88][0] ),
    .I1(\u_cpu.rf_ram.memory[89][0] ),
    .I2(\u_cpu.rf_ram.memory[90][0] ),
    .I3(\u_cpu.rf_ram.memory[91][0] ),
    .S0(_01699_),
    .S1(_01700_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06053_ (.I(_01484_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06054_ (.A1(_01698_),
    .A2(_01701_),
    .B(_01702_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06055_ (.I(_01558_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06056_ (.I(_01704_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06057_ (.I(_01616_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06058_ (.I(_01585_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06059_ (.I0(\u_cpu.rf_ram.memory[80][0] ),
    .I1(\u_cpu.rf_ram.memory[81][0] ),
    .I2(\u_cpu.rf_ram.memory[82][0] ),
    .I3(\u_cpu.rf_ram.memory[83][0] ),
    .S0(_01706_),
    .S1(_01707_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06060_ (.A1(_01705_),
    .A2(_01708_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06061_ (.I(_01466_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06062_ (.I(_01710_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06063_ (.I(_01502_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06064_ (.I(_01562_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06065_ (.I0(\u_cpu.rf_ram.memory[84][0] ),
    .I1(\u_cpu.rf_ram.memory[85][0] ),
    .I2(\u_cpu.rf_ram.memory[86][0] ),
    .I3(\u_cpu.rf_ram.memory[87][0] ),
    .S0(_01712_),
    .S1(_01713_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06066_ (.I(_01555_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06067_ (.A1(_01711_),
    .A2(_01714_),
    .B(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06068_ (.I(_01489_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06069_ (.A1(_01697_),
    .A2(_01703_),
    .B1(_01709_),
    .B2(_01716_),
    .C(_01717_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06070_ (.I(_01704_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06071_ (.I(_01540_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06072_ (.I(_01505_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06073_ (.I0(\u_cpu.rf_ram.memory[64][0] ),
    .I1(\u_cpu.rf_ram.memory[65][0] ),
    .I2(\u_cpu.rf_ram.memory[66][0] ),
    .I3(\u_cpu.rf_ram.memory[67][0] ),
    .S0(_01720_),
    .S1(_01721_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06074_ (.A1(_01719_),
    .A2(_01722_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06075_ (.I(_01710_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06076_ (.I(_01502_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06077_ (.I(_01562_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06078_ (.I0(\u_cpu.rf_ram.memory[68][0] ),
    .I1(\u_cpu.rf_ram.memory[69][0] ),
    .I2(\u_cpu.rf_ram.memory[70][0] ),
    .I3(\u_cpu.rf_ram.memory[71][0] ),
    .S0(_01725_),
    .S1(_01726_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06079_ (.I(_01555_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06080_ (.A1(_01724_),
    .A2(_01727_),
    .B(_01728_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06081_ (.I(_01704_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06082_ (.I(_01540_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06083_ (.I(_01517_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06084_ (.I0(\u_cpu.rf_ram.memory[72][0] ),
    .I1(\u_cpu.rf_ram.memory[73][0] ),
    .I2(\u_cpu.rf_ram.memory[74][0] ),
    .I3(\u_cpu.rf_ram.memory[75][0] ),
    .S0(_01731_),
    .S1(_01732_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06085_ (.A1(_01730_),
    .A2(_01733_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06086_ (.I(_01710_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06087_ (.I(_01637_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06088_ (.I0(\u_cpu.rf_ram.memory[76][0] ),
    .I1(\u_cpu.rf_ram.memory[77][0] ),
    .I2(\u_cpu.rf_ram.memory[78][0] ),
    .I3(\u_cpu.rf_ram.memory[79][0] ),
    .S0(_01515_),
    .S1(_01736_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06089_ (.I(_01484_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06090_ (.A1(_01735_),
    .A2(_01737_),
    .B(_01738_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06091_ (.I(_01577_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06092_ (.A1(_01723_),
    .A2(_01729_),
    .B1(_01734_),
    .B2(_01739_),
    .C(_01740_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06093_ (.A1(_01692_),
    .A2(_01718_),
    .A3(_01741_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06094_ (.I(_01475_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06095_ (.A1(_01691_),
    .A2(_01742_),
    .B(_01743_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06096_ (.I(_01514_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06097_ (.I(_01745_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06098_ (.I(_01746_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06099_ (.I(_01637_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06100_ (.I(_01748_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06101_ (.I0(\u_cpu.rf_ram.memory[136][0] ),
    .I1(\u_cpu.rf_ram.memory[137][0] ),
    .I2(\u_cpu.rf_ram.memory[138][0] ),
    .I3(\u_cpu.rf_ram.memory[139][0] ),
    .S0(_01747_),
    .S1(_01749_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06102_ (.A1(_01469_),
    .A2(_01750_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06103_ (.I(_01558_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06104_ (.I(_01541_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06105_ (.I(_01748_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06106_ (.I0(\u_cpu.rf_ram.memory[140][0] ),
    .I1(\u_cpu.rf_ram.memory[141][0] ),
    .I2(\u_cpu.rf_ram.memory[142][0] ),
    .I3(\u_cpu.rf_ram.memory[143][0] ),
    .S0(_01753_),
    .S1(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06107_ (.I(_01533_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06108_ (.A1(_01752_),
    .A2(_01755_),
    .B(_01756_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06109_ (.I(_01538_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06110_ (.I(_01541_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06111_ (.I(_01721_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06112_ (.I0(\u_cpu.rf_ram.memory[128][0] ),
    .I1(\u_cpu.rf_ram.memory[129][0] ),
    .I2(\u_cpu.rf_ram.memory[130][0] ),
    .I3(\u_cpu.rf_ram.memory[131][0] ),
    .S0(_01759_),
    .S1(_01760_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06113_ (.A1(_01758_),
    .A2(_01761_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06114_ (.I(_01558_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06115_ (.I(_01541_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06116_ (.I(_01721_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06117_ (.I0(\u_cpu.rf_ram.memory[132][0] ),
    .I1(\u_cpu.rf_ram.memory[133][0] ),
    .I2(\u_cpu.rf_ram.memory[134][0] ),
    .I3(\u_cpu.rf_ram.memory[135][0] ),
    .S0(_01764_),
    .S1(_01765_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06118_ (.A1(_01763_),
    .A2(_01766_),
    .B(_01574_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06119_ (.I(_01470_),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06120_ (.A1(_01751_),
    .A2(_01757_),
    .B1(_01762_),
    .B2(_01767_),
    .C(_01768_),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06121_ (.A1(_01744_),
    .A2(_01769_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06122_ (.A1(_01497_),
    .A2(_01645_),
    .B(_01770_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06123_ (.I(_01506_),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06124_ (.I0(\u_cpu.rf_ram.memory[28][1] ),
    .I1(\u_cpu.rf_ram.memory[29][1] ),
    .I2(\u_cpu.rf_ram.memory[30][1] ),
    .I3(\u_cpu.rf_ram.memory[31][1] ),
    .S0(_01504_),
    .S1(_01771_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06125_ (.A1(_01500_),
    .A2(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06126_ (.I(_01517_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06127_ (.I0(\u_cpu.rf_ram.memory[24][1] ),
    .I1(\u_cpu.rf_ram.memory[25][1] ),
    .I2(\u_cpu.rf_ram.memory[26][1] ),
    .I3(\u_cpu.rf_ram.memory[27][1] ),
    .S0(_01516_),
    .S1(_01774_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06128_ (.A1(_01513_),
    .A2(_01775_),
    .B(_01521_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06129_ (.I0(\u_cpu.rf_ram.memory[20][1] ),
    .I1(\u_cpu.rf_ram.memory[21][1] ),
    .I2(\u_cpu.rf_ram.memory[22][1] ),
    .I3(\u_cpu.rf_ram.memory[23][1] ),
    .S0(_01524_),
    .S1(_01525_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06130_ (.A1(_01523_),
    .A2(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06131_ (.I0(\u_cpu.rf_ram.memory[16][1] ),
    .I1(\u_cpu.rf_ram.memory[17][1] ),
    .I2(\u_cpu.rf_ram.memory[18][1] ),
    .I3(\u_cpu.rf_ram.memory[19][1] ),
    .S0(_01529_),
    .S1(_01530_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06132_ (.A1(_01528_),
    .A2(_01779_),
    .B(_01534_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06133_ (.A1(_01773_),
    .A2(_01776_),
    .B1(_01778_),
    .B2(_01780_),
    .C(_01490_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06134_ (.I(_01503_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06135_ (.I0(\u_cpu.rf_ram.memory[4][1] ),
    .I1(\u_cpu.rf_ram.memory[5][1] ),
    .I2(\u_cpu.rf_ram.memory[6][1] ),
    .I3(\u_cpu.rf_ram.memory[7][1] ),
    .S0(_01782_),
    .S1(_01544_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06136_ (.A1(_01539_),
    .A2(_01783_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06137_ (.I(_01512_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06138_ (.I(_01549_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06139_ (.I0(\u_cpu.rf_ram.memory[0][1] ),
    .I1(\u_cpu.rf_ram.memory[1][1] ),
    .I2(\u_cpu.rf_ram.memory[2][1] ),
    .I3(\u_cpu.rf_ram.memory[3][1] ),
    .S0(_01786_),
    .S1(_01553_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06140_ (.A1(_01785_),
    .A2(_01787_),
    .B(_01556_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06141_ (.I0(\u_cpu.rf_ram.memory[8][1] ),
    .I1(\u_cpu.rf_ram.memory[9][1] ),
    .I2(\u_cpu.rf_ram.memory[10][1] ),
    .I3(\u_cpu.rf_ram.memory[11][1] ),
    .S0(_01561_),
    .S1(_01564_),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06142_ (.A1(_01560_),
    .A2(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06143_ (.I0(\u_cpu.rf_ram.memory[12][1] ),
    .I1(\u_cpu.rf_ram.memory[13][1] ),
    .I2(\u_cpu.rf_ram.memory[14][1] ),
    .I3(\u_cpu.rf_ram.memory[15][1] ),
    .S0(_01570_),
    .S1(_01572_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06144_ (.I(_01520_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06145_ (.A1(_01567_),
    .A2(_01791_),
    .B(_01792_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06146_ (.A1(_01784_),
    .A2(_01788_),
    .B1(_01790_),
    .B2(_01793_),
    .C(_01578_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06147_ (.I(_01493_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06148_ (.I(_01628_),
    .Z(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06149_ (.I(_01583_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06150_ (.I0(\u_cpu.rf_ram.memory[36][1] ),
    .I1(\u_cpu.rf_ram.memory[37][1] ),
    .I2(\u_cpu.rf_ram.memory[38][1] ),
    .I3(\u_cpu.rf_ram.memory[39][1] ),
    .S0(_01797_),
    .S1(_01586_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06151_ (.A1(_01796_),
    .A2(_01798_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06152_ (.I0(\u_cpu.rf_ram.memory[32][1] ),
    .I1(\u_cpu.rf_ram.memory[33][1] ),
    .I2(\u_cpu.rf_ram.memory[34][1] ),
    .I3(\u_cpu.rf_ram.memory[35][1] ),
    .S0(_01590_),
    .S1(_01593_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06153_ (.I(_01532_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06154_ (.A1(_01589_),
    .A2(_01800_),
    .B(_01801_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06155_ (.I0(\u_cpu.rf_ram.memory[40][1] ),
    .I1(\u_cpu.rf_ram.memory[41][1] ),
    .I2(\u_cpu.rf_ram.memory[42][1] ),
    .I3(\u_cpu.rf_ram.memory[43][1] ),
    .S0(_01569_),
    .S1(_01601_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06156_ (.A1(_01599_),
    .A2(_01803_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06157_ (.I(_01605_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06158_ (.I0(\u_cpu.rf_ram.memory[44][1] ),
    .I1(\u_cpu.rf_ram.memory[45][1] ),
    .I2(\u_cpu.rf_ram.memory[46][1] ),
    .I3(\u_cpu.rf_ram.memory[47][1] ),
    .S0(_01805_),
    .S1(_01608_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06159_ (.I(_01610_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06160_ (.A1(_01604_),
    .A2(_01806_),
    .B(_01807_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06161_ (.A1(_01799_),
    .A2(_01802_),
    .B1(_01804_),
    .B2(_01808_),
    .C(_01613_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06162_ (.I0(\u_cpu.rf_ram.memory[60][1] ),
    .I1(\u_cpu.rf_ram.memory[61][1] ),
    .I2(\u_cpu.rf_ram.memory[62][1] ),
    .I3(\u_cpu.rf_ram.memory[63][1] ),
    .S0(_01617_),
    .S1(_01619_),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06163_ (.A1(_01615_),
    .A2(_01810_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06164_ (.I(_01592_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06165_ (.I0(\u_cpu.rf_ram.memory[56][1] ),
    .I1(\u_cpu.rf_ram.memory[57][1] ),
    .I2(\u_cpu.rf_ram.memory[58][1] ),
    .I3(\u_cpu.rf_ram.memory[59][1] ),
    .S0(_01623_),
    .S1(_01812_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06166_ (.A1(_01622_),
    .A2(_01813_),
    .B(_01626_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06167_ (.I0(\u_cpu.rf_ram.memory[52][1] ),
    .I1(\u_cpu.rf_ram.memory[53][1] ),
    .I2(\u_cpu.rf_ram.memory[54][1] ),
    .I3(\u_cpu.rf_ram.memory[55][1] ),
    .S0(_01630_),
    .S1(_01631_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06168_ (.A1(_01629_),
    .A2(_01815_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06169_ (.I0(\u_cpu.rf_ram.memory[48][1] ),
    .I1(\u_cpu.rf_ram.memory[49][1] ),
    .I2(\u_cpu.rf_ram.memory[50][1] ),
    .I3(\u_cpu.rf_ram.memory[51][1] ),
    .S0(_01636_),
    .S1(_01638_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06170_ (.A1(_01634_),
    .A2(_01817_),
    .B(_01640_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06171_ (.A1(_01811_),
    .A2(_01814_),
    .B1(_01816_),
    .B2(_01818_),
    .C(_01642_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06172_ (.A1(_01795_),
    .A2(_01809_),
    .A3(_01819_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06173_ (.A1(_01499_),
    .A2(_01781_),
    .A3(_01794_),
    .B(_01820_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06174_ (.I0(\u_cpu.rf_ram.memory[100][1] ),
    .I1(\u_cpu.rf_ram.memory[101][1] ),
    .I2(\u_cpu.rf_ram.memory[102][1] ),
    .I3(\u_cpu.rf_ram.memory[103][1] ),
    .S0(_01647_),
    .S1(_01648_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06175_ (.A1(_01646_),
    .A2(_01822_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06176_ (.I(_01592_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06177_ (.I0(\u_cpu.rf_ram.memory[96][1] ),
    .I1(\u_cpu.rf_ram.memory[97][1] ),
    .I2(\u_cpu.rf_ram.memory[98][1] ),
    .I3(\u_cpu.rf_ram.memory[99][1] ),
    .S0(_01652_),
    .S1(_01824_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06178_ (.A1(_01651_),
    .A2(_01825_),
    .B(_01654_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06179_ (.I(_01600_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06180_ (.I0(\u_cpu.rf_ram.memory[108][1] ),
    .I1(\u_cpu.rf_ram.memory[109][1] ),
    .I2(\u_cpu.rf_ram.memory[110][1] ),
    .I3(\u_cpu.rf_ram.memory[111][1] ),
    .S0(_01549_),
    .S1(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06181_ (.A1(_01656_),
    .A2(_01828_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06182_ (.I0(\u_cpu.rf_ram.memory[104][1] ),
    .I1(\u_cpu.rf_ram.memory[105][1] ),
    .I2(\u_cpu.rf_ram.memory[106][1] ),
    .I3(\u_cpu.rf_ram.memory[107][1] ),
    .S0(_01661_),
    .S1(_01571_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06183_ (.A1(_01660_),
    .A2(_01830_),
    .B(_01663_),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06184_ (.I(_01576_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06185_ (.A1(_01823_),
    .A2(_01826_),
    .B1(_01829_),
    .B2(_01831_),
    .C(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06186_ (.I0(\u_cpu.rf_ram.memory[124][1] ),
    .I1(\u_cpu.rf_ram.memory[125][1] ),
    .I2(\u_cpu.rf_ram.memory[126][1] ),
    .I3(\u_cpu.rf_ram.memory[127][1] ),
    .S0(_01668_),
    .S1(_01669_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06187_ (.A1(_01667_),
    .A2(_01834_),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06188_ (.I(_01659_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06189_ (.I(_01607_),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06190_ (.I0(\u_cpu.rf_ram.memory[120][1] ),
    .I1(\u_cpu.rf_ram.memory[121][1] ),
    .I2(\u_cpu.rf_ram.memory[122][1] ),
    .I3(\u_cpu.rf_ram.memory[123][1] ),
    .S0(_01673_),
    .S1(_01837_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06191_ (.A1(_01836_),
    .A2(_01838_),
    .B(_01676_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06192_ (.I(_01585_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06193_ (.I0(\u_cpu.rf_ram.memory[112][1] ),
    .I1(\u_cpu.rf_ram.memory[113][1] ),
    .I2(\u_cpu.rf_ram.memory[114][1] ),
    .I3(\u_cpu.rf_ram.memory[115][1] ),
    .S0(_01679_),
    .S1(_01840_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06194_ (.A1(_01678_),
    .A2(_01841_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06195_ (.I0(\u_cpu.rf_ram.memory[116][1] ),
    .I1(\u_cpu.rf_ram.memory[117][1] ),
    .I2(\u_cpu.rf_ram.memory[118][1] ),
    .I3(\u_cpu.rf_ram.memory[119][1] ),
    .S0(_01684_),
    .S1(_01685_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06196_ (.A1(_01683_),
    .A2(_01843_),
    .B(_01687_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06197_ (.A1(_01835_),
    .A2(_01839_),
    .B1(_01842_),
    .B2(_01844_),
    .C(_01689_),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06198_ (.A1(_01494_),
    .A2(_01833_),
    .A3(_01845_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06199_ (.I(_01618_),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06200_ (.I0(\u_cpu.rf_ram.memory[92][1] ),
    .I1(\u_cpu.rf_ram.memory[93][1] ),
    .I2(\u_cpu.rf_ram.memory[94][1] ),
    .I3(\u_cpu.rf_ram.memory[95][1] ),
    .S0(_01694_),
    .S1(_01847_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06201_ (.A1(_01693_),
    .A2(_01848_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06202_ (.I0(\u_cpu.rf_ram.memory[88][1] ),
    .I1(\u_cpu.rf_ram.memory[89][1] ),
    .I2(\u_cpu.rf_ram.memory[90][1] ),
    .I3(\u_cpu.rf_ram.memory[91][1] ),
    .S0(_01699_),
    .S1(_01700_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06203_ (.A1(_01698_),
    .A2(_01850_),
    .B(_01702_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06204_ (.I(_01704_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06205_ (.I0(\u_cpu.rf_ram.memory[80][1] ),
    .I1(\u_cpu.rf_ram.memory[81][1] ),
    .I2(\u_cpu.rf_ram.memory[82][1] ),
    .I3(\u_cpu.rf_ram.memory[83][1] ),
    .S0(_01706_),
    .S1(_01707_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06206_ (.A1(_01852_),
    .A2(_01853_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06207_ (.I(_01502_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06208_ (.I0(\u_cpu.rf_ram.memory[84][1] ),
    .I1(\u_cpu.rf_ram.memory[85][1] ),
    .I2(\u_cpu.rf_ram.memory[86][1] ),
    .I3(\u_cpu.rf_ram.memory[87][1] ),
    .S0(_01855_),
    .S1(_01713_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06209_ (.A1(_01711_),
    .A2(_01856_),
    .B(_01715_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06210_ (.I(_01488_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06211_ (.A1(_01849_),
    .A2(_01851_),
    .B1(_01854_),
    .B2(_01857_),
    .C(_01858_),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06212_ (.I0(\u_cpu.rf_ram.memory[64][1] ),
    .I1(\u_cpu.rf_ram.memory[65][1] ),
    .I2(\u_cpu.rf_ram.memory[66][1] ),
    .I3(\u_cpu.rf_ram.memory[67][1] ),
    .S0(_01720_),
    .S1(_01721_),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06213_ (.A1(_01719_),
    .A2(_01860_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06214_ (.I(_01710_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06215_ (.I(_01562_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06216_ (.I0(\u_cpu.rf_ram.memory[68][1] ),
    .I1(\u_cpu.rf_ram.memory[69][1] ),
    .I2(\u_cpu.rf_ram.memory[70][1] ),
    .I3(\u_cpu.rf_ram.memory[71][1] ),
    .S0(_01725_),
    .S1(_01863_),
    .Z(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06217_ (.I(_01555_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06218_ (.A1(_01862_),
    .A2(_01864_),
    .B(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06219_ (.I(_01540_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06220_ (.I0(\u_cpu.rf_ram.memory[72][1] ),
    .I1(\u_cpu.rf_ram.memory[73][1] ),
    .I2(\u_cpu.rf_ram.memory[74][1] ),
    .I3(\u_cpu.rf_ram.memory[75][1] ),
    .S0(_01867_),
    .S1(_01732_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06221_ (.A1(_01730_),
    .A2(_01868_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06222_ (.I0(\u_cpu.rf_ram.memory[76][1] ),
    .I1(\u_cpu.rf_ram.memory[77][1] ),
    .I2(\u_cpu.rf_ram.memory[78][1] ),
    .I3(\u_cpu.rf_ram.memory[79][1] ),
    .S0(_01515_),
    .S1(_01736_),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06223_ (.A1(_01735_),
    .A2(_01870_),
    .B(_01738_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06224_ (.A1(_01861_),
    .A2(_01866_),
    .B1(_01869_),
    .B2(_01871_),
    .C(_01740_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06225_ (.A1(_01692_),
    .A2(_01859_),
    .A3(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06226_ (.A1(_01846_),
    .A2(_01873_),
    .B(_01743_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06227_ (.I(_01748_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06228_ (.I0(\u_cpu.rf_ram.memory[128][1] ),
    .I1(\u_cpu.rf_ram.memory[129][1] ),
    .I2(\u_cpu.rf_ram.memory[130][1] ),
    .I3(\u_cpu.rf_ram.memory[131][1] ),
    .S0(_01747_),
    .S1(_01875_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06229_ (.A1(_01469_),
    .A2(_01876_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06230_ (.I0(\u_cpu.rf_ram.memory[132][1] ),
    .I1(\u_cpu.rf_ram.memory[133][1] ),
    .I2(\u_cpu.rf_ram.memory[134][1] ),
    .I3(\u_cpu.rf_ram.memory[135][1] ),
    .S0(_01753_),
    .S1(_01754_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06231_ (.A1(_01752_),
    .A2(_01878_),
    .B(_01485_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06232_ (.I0(\u_cpu.rf_ram.memory[136][1] ),
    .I1(\u_cpu.rf_ram.memory[137][1] ),
    .I2(\u_cpu.rf_ram.memory[138][1] ),
    .I3(\u_cpu.rf_ram.memory[139][1] ),
    .S0(_01759_),
    .S1(_01760_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06233_ (.A1(_01758_),
    .A2(_01880_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06234_ (.I0(\u_cpu.rf_ram.memory[140][1] ),
    .I1(\u_cpu.rf_ram.memory[141][1] ),
    .I2(\u_cpu.rf_ram.memory[142][1] ),
    .I3(\u_cpu.rf_ram.memory[143][1] ),
    .S0(_01764_),
    .S1(_01765_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06235_ (.A1(_01763_),
    .A2(_01882_),
    .B(_01756_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06236_ (.A1(_01877_),
    .A2(_01879_),
    .B1(_01881_),
    .B2(_01883_),
    .C(_01768_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06237_ (.A1(_01874_),
    .A2(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06238_ (.A1(_01497_),
    .A2(_01821_),
    .B(_01885_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06239_ (.I0(\u_cpu.rf_ram.memory[28][2] ),
    .I1(\u_cpu.rf_ram.memory[29][2] ),
    .I2(\u_cpu.rf_ram.memory[30][2] ),
    .I3(\u_cpu.rf_ram.memory[31][2] ),
    .S0(_01504_),
    .S1(_01771_),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06240_ (.A1(_01500_),
    .A2(_01886_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06241_ (.I0(\u_cpu.rf_ram.memory[24][2] ),
    .I1(\u_cpu.rf_ram.memory[25][2] ),
    .I2(\u_cpu.rf_ram.memory[26][2] ),
    .I3(\u_cpu.rf_ram.memory[27][2] ),
    .S0(_01516_),
    .S1(_01774_),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06242_ (.A1(_01513_),
    .A2(_01888_),
    .B(_01521_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06243_ (.I(_01467_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06244_ (.I(_01720_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06245_ (.I0(\u_cpu.rf_ram.memory[20][2] ),
    .I1(\u_cpu.rf_ram.memory[21][2] ),
    .I2(\u_cpu.rf_ram.memory[22][2] ),
    .I3(\u_cpu.rf_ram.memory[23][2] ),
    .S0(_01891_),
    .S1(_01525_),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06246_ (.A1(_01890_),
    .A2(_01892_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06247_ (.I0(\u_cpu.rf_ram.memory[16][2] ),
    .I1(\u_cpu.rf_ram.memory[17][2] ),
    .I2(\u_cpu.rf_ram.memory[18][2] ),
    .I3(\u_cpu.rf_ram.memory[19][2] ),
    .S0(_01529_),
    .S1(_01530_),
    .Z(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06248_ (.A1(_01528_),
    .A2(_01894_),
    .B(_01534_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06249_ (.A1(_01887_),
    .A2(_01889_),
    .B1(_01893_),
    .B2(_01895_),
    .C(_01490_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06250_ (.I(_01543_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06251_ (.I0(\u_cpu.rf_ram.memory[4][2] ),
    .I1(\u_cpu.rf_ram.memory[5][2] ),
    .I2(\u_cpu.rf_ram.memory[6][2] ),
    .I3(\u_cpu.rf_ram.memory[7][2] ),
    .S0(_01782_),
    .S1(_01897_),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06252_ (.A1(_01539_),
    .A2(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06253_ (.I(_01552_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06254_ (.I0(\u_cpu.rf_ram.memory[0][2] ),
    .I1(\u_cpu.rf_ram.memory[1][2] ),
    .I2(\u_cpu.rf_ram.memory[2][2] ),
    .I3(\u_cpu.rf_ram.memory[3][2] ),
    .S0(_01786_),
    .S1(_01900_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06255_ (.I(_01533_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06256_ (.A1(_01785_),
    .A2(_01901_),
    .B(_01902_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06257_ (.I0(\u_cpu.rf_ram.memory[8][2] ),
    .I1(\u_cpu.rf_ram.memory[9][2] ),
    .I2(\u_cpu.rf_ram.memory[10][2] ),
    .I3(\u_cpu.rf_ram.memory[11][2] ),
    .S0(_01561_),
    .S1(_01564_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06258_ (.A1(_01560_),
    .A2(_01904_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06259_ (.I0(\u_cpu.rf_ram.memory[12][2] ),
    .I1(\u_cpu.rf_ram.memory[13][2] ),
    .I2(\u_cpu.rf_ram.memory[14][2] ),
    .I3(\u_cpu.rf_ram.memory[15][2] ),
    .S0(_01570_),
    .S1(_01572_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06260_ (.A1(_01567_),
    .A2(_01906_),
    .B(_01792_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06261_ (.A1(_01899_),
    .A2(_01903_),
    .B1(_01905_),
    .B2(_01907_),
    .C(_01578_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06262_ (.I0(\u_cpu.rf_ram.memory[36][2] ),
    .I1(\u_cpu.rf_ram.memory[37][2] ),
    .I2(\u_cpu.rf_ram.memory[38][2] ),
    .I3(\u_cpu.rf_ram.memory[39][2] ),
    .S0(_01797_),
    .S1(_01586_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06263_ (.A1(_01796_),
    .A2(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06264_ (.I0(\u_cpu.rf_ram.memory[32][2] ),
    .I1(\u_cpu.rf_ram.memory[33][2] ),
    .I2(\u_cpu.rf_ram.memory[34][2] ),
    .I3(\u_cpu.rf_ram.memory[35][2] ),
    .S0(_01590_),
    .S1(_01593_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06265_ (.A1(_01589_),
    .A2(_01911_),
    .B(_01801_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06266_ (.I0(\u_cpu.rf_ram.memory[40][2] ),
    .I1(\u_cpu.rf_ram.memory[41][2] ),
    .I2(\u_cpu.rf_ram.memory[42][2] ),
    .I3(\u_cpu.rf_ram.memory[43][2] ),
    .S0(_01569_),
    .S1(_01601_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06267_ (.A1(_01599_),
    .A2(_01913_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06268_ (.I(_01537_),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06269_ (.I0(\u_cpu.rf_ram.memory[44][2] ),
    .I1(\u_cpu.rf_ram.memory[45][2] ),
    .I2(\u_cpu.rf_ram.memory[46][2] ),
    .I3(\u_cpu.rf_ram.memory[47][2] ),
    .S0(_01805_),
    .S1(_01608_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06270_ (.A1(_01915_),
    .A2(_01916_),
    .B(_01807_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06271_ (.A1(_01910_),
    .A2(_01912_),
    .B1(_01914_),
    .B2(_01917_),
    .C(_01613_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06272_ (.I(_01581_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06273_ (.I0(\u_cpu.rf_ram.memory[60][2] ),
    .I1(\u_cpu.rf_ram.memory[61][2] ),
    .I2(\u_cpu.rf_ram.memory[62][2] ),
    .I3(\u_cpu.rf_ram.memory[63][2] ),
    .S0(_01617_),
    .S1(_01619_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06274_ (.A1(_01919_),
    .A2(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06275_ (.I0(\u_cpu.rf_ram.memory[56][2] ),
    .I1(\u_cpu.rf_ram.memory[57][2] ),
    .I2(\u_cpu.rf_ram.memory[58][2] ),
    .I3(\u_cpu.rf_ram.memory[59][2] ),
    .S0(_01623_),
    .S1(_01812_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06276_ (.A1(_01622_),
    .A2(_01922_),
    .B(_01626_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06277_ (.I0(\u_cpu.rf_ram.memory[52][2] ),
    .I1(\u_cpu.rf_ram.memory[53][2] ),
    .I2(\u_cpu.rf_ram.memory[54][2] ),
    .I3(\u_cpu.rf_ram.memory[55][2] ),
    .S0(_01630_),
    .S1(_01631_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06278_ (.A1(_01629_),
    .A2(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06279_ (.I(_01598_),
    .Z(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06280_ (.I(_01637_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06281_ (.I0(\u_cpu.rf_ram.memory[48][2] ),
    .I1(\u_cpu.rf_ram.memory[49][2] ),
    .I2(\u_cpu.rf_ram.memory[50][2] ),
    .I3(\u_cpu.rf_ram.memory[51][2] ),
    .S0(_01636_),
    .S1(_01927_),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06282_ (.I(_01595_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06283_ (.A1(_01926_),
    .A2(_01928_),
    .B(_01929_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06284_ (.A1(_01921_),
    .A2(_01923_),
    .B1(_01925_),
    .B2(_01930_),
    .C(_01642_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06285_ (.A1(_01795_),
    .A2(_01918_),
    .A3(_01931_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06286_ (.A1(_01499_),
    .A2(_01896_),
    .A3(_01908_),
    .B(_01932_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06287_ (.I(_01568_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06288_ (.I0(\u_cpu.rf_ram.memory[100][2] ),
    .I1(\u_cpu.rf_ram.memory[101][2] ),
    .I2(\u_cpu.rf_ram.memory[102][2] ),
    .I3(\u_cpu.rf_ram.memory[103][2] ),
    .S0(_01934_),
    .S1(_01648_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06289_ (.A1(_01646_),
    .A2(_01935_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06290_ (.I(_01511_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06291_ (.I(_01548_),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06292_ (.I0(\u_cpu.rf_ram.memory[96][2] ),
    .I1(\u_cpu.rf_ram.memory[97][2] ),
    .I2(\u_cpu.rf_ram.memory[98][2] ),
    .I3(\u_cpu.rf_ram.memory[99][2] ),
    .S0(_01938_),
    .S1(_01824_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06293_ (.A1(_01937_),
    .A2(_01939_),
    .B(_01654_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06294_ (.I(_01710_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06295_ (.I0(\u_cpu.rf_ram.memory[108][2] ),
    .I1(\u_cpu.rf_ram.memory[109][2] ),
    .I2(\u_cpu.rf_ram.memory[110][2] ),
    .I3(\u_cpu.rf_ram.memory[111][2] ),
    .S0(_01549_),
    .S1(_01827_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06296_ (.A1(_01941_),
    .A2(_01942_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06297_ (.I0(\u_cpu.rf_ram.memory[104][2] ),
    .I1(\u_cpu.rf_ram.memory[105][2] ),
    .I2(\u_cpu.rf_ram.memory[106][2] ),
    .I3(\u_cpu.rf_ram.memory[107][2] ),
    .S0(_01661_),
    .S1(_01571_),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06298_ (.A1(_01660_),
    .A2(_01944_),
    .B(_01663_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06299_ (.A1(_01936_),
    .A2(_01940_),
    .B1(_01943_),
    .B2(_01945_),
    .C(_01832_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06300_ (.I(_01616_),
    .Z(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06301_ (.I0(\u_cpu.rf_ram.memory[124][2] ),
    .I1(\u_cpu.rf_ram.memory[125][2] ),
    .I2(\u_cpu.rf_ram.memory[126][2] ),
    .I3(\u_cpu.rf_ram.memory[127][2] ),
    .S0(_01947_),
    .S1(_01669_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06302_ (.A1(_01667_),
    .A2(_01948_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06303_ (.I0(\u_cpu.rf_ram.memory[120][2] ),
    .I1(\u_cpu.rf_ram.memory[121][2] ),
    .I2(\u_cpu.rf_ram.memory[122][2] ),
    .I3(\u_cpu.rf_ram.memory[123][2] ),
    .S0(_01673_),
    .S1(_01837_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06304_ (.A1(_01836_),
    .A2(_01950_),
    .B(_01676_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06305_ (.I0(\u_cpu.rf_ram.memory[112][2] ),
    .I1(\u_cpu.rf_ram.memory[113][2] ),
    .I2(\u_cpu.rf_ram.memory[114][2] ),
    .I3(\u_cpu.rf_ram.memory[115][2] ),
    .S0(_01679_),
    .S1(_01840_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06306_ (.A1(_01678_),
    .A2(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06307_ (.I0(\u_cpu.rf_ram.memory[116][2] ),
    .I1(\u_cpu.rf_ram.memory[117][2] ),
    .I2(\u_cpu.rf_ram.memory[118][2] ),
    .I3(\u_cpu.rf_ram.memory[119][2] ),
    .S0(_01684_),
    .S1(_01685_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06308_ (.A1(_01683_),
    .A2(_01954_),
    .B(_01687_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06309_ (.A1(_01949_),
    .A2(_01951_),
    .B1(_01953_),
    .B2(_01955_),
    .C(_01689_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06310_ (.A1(_01494_),
    .A2(_01946_),
    .A3(_01956_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06311_ (.I(_01498_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06312_ (.I0(\u_cpu.rf_ram.memory[92][2] ),
    .I1(\u_cpu.rf_ram.memory[93][2] ),
    .I2(\u_cpu.rf_ram.memory[94][2] ),
    .I3(\u_cpu.rf_ram.memory[95][2] ),
    .S0(_01694_),
    .S1(_01847_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06313_ (.A1(_01693_),
    .A2(_01959_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06314_ (.I(_01635_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06315_ (.I0(\u_cpu.rf_ram.memory[88][2] ),
    .I1(\u_cpu.rf_ram.memory[89][2] ),
    .I2(\u_cpu.rf_ram.memory[90][2] ),
    .I3(\u_cpu.rf_ram.memory[91][2] ),
    .S0(_01961_),
    .S1(_01700_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06316_ (.I(_01610_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06317_ (.A1(_01698_),
    .A2(_01962_),
    .B(_01963_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06318_ (.I(_01585_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06319_ (.I0(\u_cpu.rf_ram.memory[80][2] ),
    .I1(\u_cpu.rf_ram.memory[81][2] ),
    .I2(\u_cpu.rf_ram.memory[82][2] ),
    .I3(\u_cpu.rf_ram.memory[83][2] ),
    .S0(_01706_),
    .S1(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06320_ (.A1(_01852_),
    .A2(_01966_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06321_ (.I0(\u_cpu.rf_ram.memory[84][2] ),
    .I1(\u_cpu.rf_ram.memory[85][2] ),
    .I2(\u_cpu.rf_ram.memory[86][2] ),
    .I3(\u_cpu.rf_ram.memory[87][2] ),
    .S0(_01855_),
    .S1(_01713_),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06322_ (.A1(_01711_),
    .A2(_01968_),
    .B(_01715_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06323_ (.A1(_01960_),
    .A2(_01964_),
    .B1(_01967_),
    .B2(_01969_),
    .C(_01858_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06324_ (.I(_01704_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06325_ (.I(_01517_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06326_ (.I0(\u_cpu.rf_ram.memory[64][2] ),
    .I1(\u_cpu.rf_ram.memory[65][2] ),
    .I2(\u_cpu.rf_ram.memory[66][2] ),
    .I3(\u_cpu.rf_ram.memory[67][2] ),
    .S0(_01720_),
    .S1(_01972_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06327_ (.A1(_01971_),
    .A2(_01973_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06328_ (.I0(\u_cpu.rf_ram.memory[68][2] ),
    .I1(\u_cpu.rf_ram.memory[69][2] ),
    .I2(\u_cpu.rf_ram.memory[70][2] ),
    .I3(\u_cpu.rf_ram.memory[71][2] ),
    .S0(_01725_),
    .S1(_01863_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06329_ (.A1(_01862_),
    .A2(_01975_),
    .B(_01865_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06330_ (.I0(\u_cpu.rf_ram.memory[72][2] ),
    .I1(\u_cpu.rf_ram.memory[73][2] ),
    .I2(\u_cpu.rf_ram.memory[74][2] ),
    .I3(\u_cpu.rf_ram.memory[75][2] ),
    .S0(_01867_),
    .S1(_01732_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06331_ (.A1(_01730_),
    .A2(_01977_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06332_ (.I(_01502_),
    .Z(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06333_ (.I0(\u_cpu.rf_ram.memory[76][2] ),
    .I1(\u_cpu.rf_ram.memory[77][2] ),
    .I2(\u_cpu.rf_ram.memory[78][2] ),
    .I3(\u_cpu.rf_ram.memory[79][2] ),
    .S0(_01979_),
    .S1(_01736_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06334_ (.A1(_01735_),
    .A2(_01980_),
    .B(_01738_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06335_ (.I(_01577_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06336_ (.A1(_01974_),
    .A2(_01976_),
    .B1(_01978_),
    .B2(_01981_),
    .C(_01982_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06337_ (.A1(_01958_),
    .A2(_01970_),
    .A3(_01983_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06338_ (.A1(_01957_),
    .A2(_01984_),
    .B(_01743_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06339_ (.I0(\u_cpu.rf_ram.memory[136][2] ),
    .I1(\u_cpu.rf_ram.memory[137][2] ),
    .I2(\u_cpu.rf_ram.memory[138][2] ),
    .I3(\u_cpu.rf_ram.memory[139][2] ),
    .S0(_01747_),
    .S1(_01875_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06340_ (.A1(_01469_),
    .A2(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06341_ (.I0(\u_cpu.rf_ram.memory[140][2] ),
    .I1(\u_cpu.rf_ram.memory[141][2] ),
    .I2(\u_cpu.rf_ram.memory[142][2] ),
    .I3(\u_cpu.rf_ram.memory[143][2] ),
    .S0(_01753_),
    .S1(_01754_),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06342_ (.A1(_01752_),
    .A2(_01988_),
    .B(_01756_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06343_ (.I0(\u_cpu.rf_ram.memory[128][2] ),
    .I1(\u_cpu.rf_ram.memory[129][2] ),
    .I2(\u_cpu.rf_ram.memory[130][2] ),
    .I3(\u_cpu.rf_ram.memory[131][2] ),
    .S0(_01759_),
    .S1(_01760_),
    .Z(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06344_ (.A1(_01758_),
    .A2(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06345_ (.I(_01558_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06346_ (.I(_01541_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06347_ (.I0(\u_cpu.rf_ram.memory[132][2] ),
    .I1(\u_cpu.rf_ram.memory[133][2] ),
    .I2(\u_cpu.rf_ram.memory[134][2] ),
    .I3(\u_cpu.rf_ram.memory[135][2] ),
    .S0(_01993_),
    .S1(_01765_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06348_ (.A1(_01992_),
    .A2(_01994_),
    .B(_01574_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06349_ (.A1(_01987_),
    .A2(_01989_),
    .B1(_01991_),
    .B2(_01995_),
    .C(_01768_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06350_ (.A1(_01985_),
    .A2(_01996_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06351_ (.A1(_01497_),
    .A2(_01933_),
    .B(_01997_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06352_ (.I0(\u_cpu.rf_ram.memory[28][3] ),
    .I1(\u_cpu.rf_ram.memory[29][3] ),
    .I2(\u_cpu.rf_ram.memory[30][3] ),
    .I3(\u_cpu.rf_ram.memory[31][3] ),
    .S0(_01504_),
    .S1(_01771_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06353_ (.A1(_01500_),
    .A2(_01998_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06354_ (.I0(\u_cpu.rf_ram.memory[24][3] ),
    .I1(\u_cpu.rf_ram.memory[25][3] ),
    .I2(\u_cpu.rf_ram.memory[26][3] ),
    .I3(\u_cpu.rf_ram.memory[27][3] ),
    .S0(_01516_),
    .S1(_01774_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06355_ (.I(_01484_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06356_ (.A1(_01513_),
    .A2(_02000_),
    .B(_02001_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06357_ (.I(_01736_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06358_ (.I0(\u_cpu.rf_ram.memory[20][3] ),
    .I1(\u_cpu.rf_ram.memory[21][3] ),
    .I2(\u_cpu.rf_ram.memory[22][3] ),
    .I3(\u_cpu.rf_ram.memory[23][3] ),
    .S0(_01891_),
    .S1(_02003_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06359_ (.A1(_01890_),
    .A2(_02004_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06360_ (.I(_01512_),
    .Z(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06361_ (.I(_01515_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06362_ (.I0(\u_cpu.rf_ram.memory[16][3] ),
    .I1(\u_cpu.rf_ram.memory[17][3] ),
    .I2(\u_cpu.rf_ram.memory[18][3] ),
    .I3(\u_cpu.rf_ram.memory[19][3] ),
    .S0(_02007_),
    .S1(_01530_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06363_ (.A1(_02006_),
    .A2(_02008_),
    .B(_01534_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06364_ (.A1(_01999_),
    .A2(_02002_),
    .B1(_02005_),
    .B2(_02009_),
    .C(_01490_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06365_ (.I(_01538_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06366_ (.I0(\u_cpu.rf_ram.memory[4][3] ),
    .I1(\u_cpu.rf_ram.memory[5][3] ),
    .I2(\u_cpu.rf_ram.memory[6][3] ),
    .I3(\u_cpu.rf_ram.memory[7][3] ),
    .S0(_01782_),
    .S1(_01897_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06367_ (.A1(_02011_),
    .A2(_02012_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06368_ (.I0(\u_cpu.rf_ram.memory[0][3] ),
    .I1(\u_cpu.rf_ram.memory[1][3] ),
    .I2(\u_cpu.rf_ram.memory[2][3] ),
    .I3(\u_cpu.rf_ram.memory[3][3] ),
    .S0(_01786_),
    .S1(_01900_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06369_ (.A1(_01785_),
    .A2(_02014_),
    .B(_01902_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06370_ (.I(_01503_),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06371_ (.I0(\u_cpu.rf_ram.memory[8][3] ),
    .I1(\u_cpu.rf_ram.memory[9][3] ),
    .I2(\u_cpu.rf_ram.memory[10][3] ),
    .I3(\u_cpu.rf_ram.memory[11][3] ),
    .S0(_02016_),
    .S1(_01564_),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06372_ (.A1(_01560_),
    .A2(_02017_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06373_ (.I0(\u_cpu.rf_ram.memory[12][3] ),
    .I1(\u_cpu.rf_ram.memory[13][3] ),
    .I2(\u_cpu.rf_ram.memory[14][3] ),
    .I3(\u_cpu.rf_ram.memory[15][3] ),
    .S0(_01570_),
    .S1(_01572_),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06374_ (.A1(_01567_),
    .A2(_02019_),
    .B(_01792_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06375_ (.A1(_02013_),
    .A2(_02015_),
    .B1(_02018_),
    .B2(_02020_),
    .C(_01578_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06376_ (.I0(\u_cpu.rf_ram.memory[36][3] ),
    .I1(\u_cpu.rf_ram.memory[37][3] ),
    .I2(\u_cpu.rf_ram.memory[38][3] ),
    .I3(\u_cpu.rf_ram.memory[39][3] ),
    .S0(_01797_),
    .S1(_01586_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06377_ (.A1(_01796_),
    .A2(_02022_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06378_ (.I(_01592_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06379_ (.I0(\u_cpu.rf_ram.memory[32][3] ),
    .I1(\u_cpu.rf_ram.memory[33][3] ),
    .I2(\u_cpu.rf_ram.memory[34][3] ),
    .I3(\u_cpu.rf_ram.memory[35][3] ),
    .S0(_01590_),
    .S1(_02024_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06380_ (.A1(_01589_),
    .A2(_02025_),
    .B(_01801_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06381_ (.I(_01568_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06382_ (.I0(\u_cpu.rf_ram.memory[40][3] ),
    .I1(\u_cpu.rf_ram.memory[41][3] ),
    .I2(\u_cpu.rf_ram.memory[42][3] ),
    .I3(\u_cpu.rf_ram.memory[43][3] ),
    .S0(_02027_),
    .S1(_01601_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06383_ (.A1(_01599_),
    .A2(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06384_ (.I(_01607_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06385_ (.I0(\u_cpu.rf_ram.memory[44][3] ),
    .I1(\u_cpu.rf_ram.memory[45][3] ),
    .I2(\u_cpu.rf_ram.memory[46][3] ),
    .I3(\u_cpu.rf_ram.memory[47][3] ),
    .S0(_01805_),
    .S1(_02030_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06386_ (.A1(_01915_),
    .A2(_02031_),
    .B(_01807_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06387_ (.A1(_02023_),
    .A2(_02026_),
    .B1(_02029_),
    .B2(_02032_),
    .C(_01613_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06388_ (.I(_01618_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06389_ (.I0(\u_cpu.rf_ram.memory[60][3] ),
    .I1(\u_cpu.rf_ram.memory[61][3] ),
    .I2(\u_cpu.rf_ram.memory[62][3] ),
    .I3(\u_cpu.rf_ram.memory[63][3] ),
    .S0(_01617_),
    .S1(_02034_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06390_ (.A1(_01919_),
    .A2(_02035_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06391_ (.I0(\u_cpu.rf_ram.memory[56][3] ),
    .I1(\u_cpu.rf_ram.memory[57][3] ),
    .I2(\u_cpu.rf_ram.memory[58][3] ),
    .I3(\u_cpu.rf_ram.memory[59][3] ),
    .S0(_01623_),
    .S1(_01812_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06392_ (.A1(_01622_),
    .A2(_02037_),
    .B(_01626_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06393_ (.I(_01628_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06394_ (.I(_01600_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06395_ (.I0(\u_cpu.rf_ram.memory[52][3] ),
    .I1(\u_cpu.rf_ram.memory[53][3] ),
    .I2(\u_cpu.rf_ram.memory[54][3] ),
    .I3(\u_cpu.rf_ram.memory[55][3] ),
    .S0(_01630_),
    .S1(_02040_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06396_ (.A1(_02039_),
    .A2(_02041_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06397_ (.I0(\u_cpu.rf_ram.memory[48][3] ),
    .I1(\u_cpu.rf_ram.memory[49][3] ),
    .I2(\u_cpu.rf_ram.memory[50][3] ),
    .I3(\u_cpu.rf_ram.memory[51][3] ),
    .S0(_01636_),
    .S1(_01927_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06398_ (.A1(_01926_),
    .A2(_02043_),
    .B(_01929_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06399_ (.A1(_02036_),
    .A2(_02038_),
    .B1(_02042_),
    .B2(_02044_),
    .C(_01642_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06400_ (.A1(_01795_),
    .A2(_02033_),
    .A3(_02045_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06401_ (.A1(_01499_),
    .A2(_02010_),
    .A3(_02021_),
    .B(_02046_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06402_ (.I0(\u_cpu.rf_ram.memory[100][3] ),
    .I1(\u_cpu.rf_ram.memory[101][3] ),
    .I2(\u_cpu.rf_ram.memory[102][3] ),
    .I3(\u_cpu.rf_ram.memory[103][3] ),
    .S0(_01934_),
    .S1(_01648_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06403_ (.A1(_01646_),
    .A2(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06404_ (.I0(\u_cpu.rf_ram.memory[96][3] ),
    .I1(\u_cpu.rf_ram.memory[97][3] ),
    .I2(\u_cpu.rf_ram.memory[98][3] ),
    .I3(\u_cpu.rf_ram.memory[99][3] ),
    .S0(_01938_),
    .S1(_01824_),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06405_ (.A1(_01937_),
    .A2(_02050_),
    .B(_01654_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06406_ (.I(_01568_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06407_ (.I0(\u_cpu.rf_ram.memory[108][3] ),
    .I1(\u_cpu.rf_ram.memory[109][3] ),
    .I2(\u_cpu.rf_ram.memory[110][3] ),
    .I3(\u_cpu.rf_ram.memory[111][3] ),
    .S0(_02052_),
    .S1(_01827_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06408_ (.A1(_01941_),
    .A2(_02053_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06409_ (.I(_01659_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06410_ (.I(_01605_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06411_ (.I0(\u_cpu.rf_ram.memory[104][3] ),
    .I1(\u_cpu.rf_ram.memory[105][3] ),
    .I2(\u_cpu.rf_ram.memory[106][3] ),
    .I3(\u_cpu.rf_ram.memory[107][3] ),
    .S0(_02056_),
    .S1(_01571_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06412_ (.I(_01483_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06413_ (.A1(_02055_),
    .A2(_02057_),
    .B(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06414_ (.A1(_02049_),
    .A2(_02051_),
    .B1(_02054_),
    .B2(_02059_),
    .C(_01832_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06415_ (.I0(\u_cpu.rf_ram.memory[124][3] ),
    .I1(\u_cpu.rf_ram.memory[125][3] ),
    .I2(\u_cpu.rf_ram.memory[126][3] ),
    .I3(\u_cpu.rf_ram.memory[127][3] ),
    .S0(_01947_),
    .S1(_01669_),
    .Z(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06416_ (.A1(_01667_),
    .A2(_02061_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06417_ (.I0(\u_cpu.rf_ram.memory[120][3] ),
    .I1(\u_cpu.rf_ram.memory[121][3] ),
    .I2(\u_cpu.rf_ram.memory[122][3] ),
    .I3(\u_cpu.rf_ram.memory[123][3] ),
    .S0(_01673_),
    .S1(_01837_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06418_ (.A1(_01836_),
    .A2(_02063_),
    .B(_01676_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06419_ (.I(_01598_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06420_ (.I(_01583_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06421_ (.I0(\u_cpu.rf_ram.memory[112][3] ),
    .I1(\u_cpu.rf_ram.memory[113][3] ),
    .I2(\u_cpu.rf_ram.memory[114][3] ),
    .I3(\u_cpu.rf_ram.memory[115][3] ),
    .S0(_02066_),
    .S1(_01840_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06422_ (.A1(_02065_),
    .A2(_02067_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06423_ (.I(_01635_),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06424_ (.I0(\u_cpu.rf_ram.memory[116][3] ),
    .I1(\u_cpu.rf_ram.memory[117][3] ),
    .I2(\u_cpu.rf_ram.memory[118][3] ),
    .I3(\u_cpu.rf_ram.memory[119][3] ),
    .S0(_02069_),
    .S1(_01685_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06425_ (.A1(_01683_),
    .A2(_02070_),
    .B(_01687_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06426_ (.I(_01488_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06427_ (.A1(_02062_),
    .A2(_02064_),
    .B1(_02068_),
    .B2(_02071_),
    .C(_02072_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06428_ (.A1(_01494_),
    .A2(_02060_),
    .A3(_02073_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06429_ (.I(_01616_),
    .Z(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06430_ (.I0(\u_cpu.rf_ram.memory[92][3] ),
    .I1(\u_cpu.rf_ram.memory[93][3] ),
    .I2(\u_cpu.rf_ram.memory[94][3] ),
    .I3(\u_cpu.rf_ram.memory[95][3] ),
    .S0(_02075_),
    .S1(_01847_),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06431_ (.A1(_01693_),
    .A2(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06432_ (.I0(\u_cpu.rf_ram.memory[88][3] ),
    .I1(\u_cpu.rf_ram.memory[89][3] ),
    .I2(\u_cpu.rf_ram.memory[90][3] ),
    .I3(\u_cpu.rf_ram.memory[91][3] ),
    .S0(_01961_),
    .S1(_01700_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06433_ (.A1(_01698_),
    .A2(_02078_),
    .B(_01963_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06434_ (.I0(\u_cpu.rf_ram.memory[80][3] ),
    .I1(\u_cpu.rf_ram.memory[81][3] ),
    .I2(\u_cpu.rf_ram.memory[82][3] ),
    .I3(\u_cpu.rf_ram.memory[83][3] ),
    .S0(_01706_),
    .S1(_01965_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06435_ (.A1(_01852_),
    .A2(_02080_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06436_ (.I(_01537_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06437_ (.I(_01562_),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06438_ (.I0(\u_cpu.rf_ram.memory[84][3] ),
    .I1(\u_cpu.rf_ram.memory[85][3] ),
    .I2(\u_cpu.rf_ram.memory[86][3] ),
    .I3(\u_cpu.rf_ram.memory[87][3] ),
    .S0(_01855_),
    .S1(_02083_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06439_ (.I(_01555_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06440_ (.A1(_02082_),
    .A2(_02084_),
    .B(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06441_ (.A1(_02077_),
    .A2(_02079_),
    .B1(_02081_),
    .B2(_02086_),
    .C(_01858_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06442_ (.I0(\u_cpu.rf_ram.memory[64][3] ),
    .I1(\u_cpu.rf_ram.memory[65][3] ),
    .I2(\u_cpu.rf_ram.memory[66][3] ),
    .I3(\u_cpu.rf_ram.memory[67][3] ),
    .S0(_01720_),
    .S1(_01972_),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06443_ (.A1(_01971_),
    .A2(_02088_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06444_ (.I0(\u_cpu.rf_ram.memory[68][3] ),
    .I1(\u_cpu.rf_ram.memory[69][3] ),
    .I2(\u_cpu.rf_ram.memory[70][3] ),
    .I3(\u_cpu.rf_ram.memory[71][3] ),
    .S0(_01725_),
    .S1(_01863_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06445_ (.A1(_01862_),
    .A2(_02090_),
    .B(_01865_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06446_ (.I0(\u_cpu.rf_ram.memory[72][3] ),
    .I1(\u_cpu.rf_ram.memory[73][3] ),
    .I2(\u_cpu.rf_ram.memory[74][3] ),
    .I3(\u_cpu.rf_ram.memory[75][3] ),
    .S0(_01867_),
    .S1(_01732_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06447_ (.A1(_01730_),
    .A2(_02092_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06448_ (.I0(\u_cpu.rf_ram.memory[76][3] ),
    .I1(\u_cpu.rf_ram.memory[77][3] ),
    .I2(\u_cpu.rf_ram.memory[78][3] ),
    .I3(\u_cpu.rf_ram.memory[79][3] ),
    .S0(_01979_),
    .S1(_01736_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06449_ (.A1(_01735_),
    .A2(_02094_),
    .B(_01738_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06450_ (.A1(_02089_),
    .A2(_02091_),
    .B1(_02093_),
    .B2(_02095_),
    .C(_01982_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06451_ (.A1(_01958_),
    .A2(_02087_),
    .A3(_02096_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06452_ (.A1(_02074_),
    .A2(_02097_),
    .B(_01743_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06453_ (.I0(\u_cpu.rf_ram.memory[128][3] ),
    .I1(\u_cpu.rf_ram.memory[129][3] ),
    .I2(\u_cpu.rf_ram.memory[130][3] ),
    .I3(\u_cpu.rf_ram.memory[131][3] ),
    .S0(_01747_),
    .S1(_01875_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06454_ (.A1(_01469_),
    .A2(_02099_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06455_ (.I(_01746_),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06456_ (.I0(\u_cpu.rf_ram.memory[132][3] ),
    .I1(\u_cpu.rf_ram.memory[133][3] ),
    .I2(\u_cpu.rf_ram.memory[134][3] ),
    .I3(\u_cpu.rf_ram.memory[135][3] ),
    .S0(_02101_),
    .S1(_01754_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06457_ (.A1(_01752_),
    .A2(_02102_),
    .B(_01485_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06458_ (.I0(\u_cpu.rf_ram.memory[136][3] ),
    .I1(\u_cpu.rf_ram.memory[137][3] ),
    .I2(\u_cpu.rf_ram.memory[138][3] ),
    .I3(\u_cpu.rf_ram.memory[139][3] ),
    .S0(_01759_),
    .S1(_01760_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06459_ (.A1(_01758_),
    .A2(_02104_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06460_ (.I(_01721_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06461_ (.I0(\u_cpu.rf_ram.memory[140][3] ),
    .I1(\u_cpu.rf_ram.memory[141][3] ),
    .I2(\u_cpu.rf_ram.memory[142][3] ),
    .I3(\u_cpu.rf_ram.memory[143][3] ),
    .S0(_01993_),
    .S1(_02106_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06462_ (.A1(_01992_),
    .A2(_02107_),
    .B(_01556_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06463_ (.A1(_02100_),
    .A2(_02103_),
    .B1(_02105_),
    .B2(_02108_),
    .C(_01768_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06464_ (.A1(_02098_),
    .A2(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06465_ (.A1(_01497_),
    .A2(_02047_),
    .B(_02110_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06466_ (.I0(\u_cpu.rf_ram.memory[28][4] ),
    .I1(\u_cpu.rf_ram.memory[29][4] ),
    .I2(\u_cpu.rf_ram.memory[30][4] ),
    .I3(\u_cpu.rf_ram.memory[31][4] ),
    .S0(_01504_),
    .S1(_01771_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06467_ (.A1(_01500_),
    .A2(_02111_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06468_ (.I0(\u_cpu.rf_ram.memory[24][4] ),
    .I1(\u_cpu.rf_ram.memory[25][4] ),
    .I2(\u_cpu.rf_ram.memory[26][4] ),
    .I3(\u_cpu.rf_ram.memory[27][4] ),
    .S0(_01516_),
    .S1(_01774_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06469_ (.A1(_01513_),
    .A2(_02113_),
    .B(_02001_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06470_ (.I0(\u_cpu.rf_ram.memory[20][4] ),
    .I1(\u_cpu.rf_ram.memory[21][4] ),
    .I2(\u_cpu.rf_ram.memory[22][4] ),
    .I3(\u_cpu.rf_ram.memory[23][4] ),
    .S0(_01891_),
    .S1(_02003_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06471_ (.A1(_01890_),
    .A2(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06472_ (.I0(\u_cpu.rf_ram.memory[16][4] ),
    .I1(\u_cpu.rf_ram.memory[17][4] ),
    .I2(\u_cpu.rf_ram.memory[18][4] ),
    .I3(\u_cpu.rf_ram.memory[19][4] ),
    .S0(_02007_),
    .S1(_01518_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06473_ (.A1(_02006_),
    .A2(_02117_),
    .B(_01728_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06474_ (.A1(_02112_),
    .A2(_02114_),
    .B1(_02116_),
    .B2(_02118_),
    .C(_01717_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06475_ (.I0(\u_cpu.rf_ram.memory[4][4] ),
    .I1(\u_cpu.rf_ram.memory[5][4] ),
    .I2(\u_cpu.rf_ram.memory[6][4] ),
    .I3(\u_cpu.rf_ram.memory[7][4] ),
    .S0(_01782_),
    .S1(_01897_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06476_ (.A1(_02011_),
    .A2(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06477_ (.I0(\u_cpu.rf_ram.memory[0][4] ),
    .I1(\u_cpu.rf_ram.memory[1][4] ),
    .I2(\u_cpu.rf_ram.memory[2][4] ),
    .I3(\u_cpu.rf_ram.memory[3][4] ),
    .S0(_01786_),
    .S1(_01900_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06478_ (.A1(_01785_),
    .A2(_02122_),
    .B(_01902_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06479_ (.I0(\u_cpu.rf_ram.memory[8][4] ),
    .I1(\u_cpu.rf_ram.memory[9][4] ),
    .I2(\u_cpu.rf_ram.memory[10][4] ),
    .I3(\u_cpu.rf_ram.memory[11][4] ),
    .S0(_02016_),
    .S1(_01507_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06480_ (.A1(_01547_),
    .A2(_02124_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06481_ (.I0(\u_cpu.rf_ram.memory[12][4] ),
    .I1(\u_cpu.rf_ram.memory[13][4] ),
    .I2(\u_cpu.rf_ram.memory[14][4] ),
    .I3(\u_cpu.rf_ram.memory[15][4] ),
    .S0(_01550_),
    .S1(_01572_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06482_ (.A1(_01468_),
    .A2(_02126_),
    .B(_01792_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06483_ (.A1(_02121_),
    .A2(_02123_),
    .B1(_02125_),
    .B2(_02127_),
    .C(_01578_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06484_ (.I0(\u_cpu.rf_ram.memory[36][4] ),
    .I1(\u_cpu.rf_ram.memory[37][4] ),
    .I2(\u_cpu.rf_ram.memory[38][4] ),
    .I3(\u_cpu.rf_ram.memory[39][4] ),
    .S0(_01797_),
    .S1(_01680_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06485_ (.A1(_01796_),
    .A2(_02129_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06486_ (.I0(\u_cpu.rf_ram.memory[32][4] ),
    .I1(\u_cpu.rf_ram.memory[33][4] ),
    .I2(\u_cpu.rf_ram.memory[34][4] ),
    .I3(\u_cpu.rf_ram.memory[35][4] ),
    .S0(_01745_),
    .S1(_02024_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06487_ (.A1(_01559_),
    .A2(_02131_),
    .B(_01801_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06488_ (.I0(\u_cpu.rf_ram.memory[40][4] ),
    .I1(\u_cpu.rf_ram.memory[41][4] ),
    .I2(\u_cpu.rf_ram.memory[42][4] ),
    .I3(\u_cpu.rf_ram.memory[43][4] ),
    .S0(_02027_),
    .S1(_01601_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06489_ (.A1(_01599_),
    .A2(_02133_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06490_ (.I0(\u_cpu.rf_ram.memory[44][4] ),
    .I1(\u_cpu.rf_ram.memory[45][4] ),
    .I2(\u_cpu.rf_ram.memory[46][4] ),
    .I3(\u_cpu.rf_ram.memory[47][4] ),
    .S0(_01805_),
    .S1(_02030_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06491_ (.A1(_01915_),
    .A2(_02135_),
    .B(_01807_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06492_ (.A1(_02130_),
    .A2(_02132_),
    .B1(_02134_),
    .B2(_02136_),
    .C(_01665_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06493_ (.I0(\u_cpu.rf_ram.memory[60][4] ),
    .I1(\u_cpu.rf_ram.memory[61][4] ),
    .I2(\u_cpu.rf_ram.memory[62][4] ),
    .I3(\u_cpu.rf_ram.memory[63][4] ),
    .S0(_01617_),
    .S1(_02034_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06494_ (.A1(_01919_),
    .A2(_02138_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06495_ (.I0(\u_cpu.rf_ram.memory[56][4] ),
    .I1(\u_cpu.rf_ram.memory[57][4] ),
    .I2(\u_cpu.rf_ram.memory[58][4] ),
    .I3(\u_cpu.rf_ram.memory[59][4] ),
    .S0(_01623_),
    .S1(_01812_),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06496_ (.A1(_01622_),
    .A2(_02140_),
    .B(_01626_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06497_ (.I0(\u_cpu.rf_ram.memory[52][4] ),
    .I1(\u_cpu.rf_ram.memory[53][4] ),
    .I2(\u_cpu.rf_ram.memory[54][4] ),
    .I3(\u_cpu.rf_ram.memory[55][4] ),
    .S0(_01630_),
    .S1(_02040_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06498_ (.A1(_02039_),
    .A2(_02142_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06499_ (.I0(\u_cpu.rf_ram.memory[48][4] ),
    .I1(\u_cpu.rf_ram.memory[49][4] ),
    .I2(\u_cpu.rf_ram.memory[50][4] ),
    .I3(\u_cpu.rf_ram.memory[51][4] ),
    .S0(_01636_),
    .S1(_01927_),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06500_ (.A1(_01926_),
    .A2(_02144_),
    .B(_01929_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06501_ (.A1(_02139_),
    .A2(_02141_),
    .B1(_02143_),
    .B2(_02145_),
    .C(_01642_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06502_ (.A1(_01795_),
    .A2(_02137_),
    .A3(_02146_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06503_ (.A1(_01499_),
    .A2(_02119_),
    .A3(_02128_),
    .B(_02147_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06504_ (.I0(\u_cpu.rf_ram.memory[100][4] ),
    .I1(\u_cpu.rf_ram.memory[101][4] ),
    .I2(\u_cpu.rf_ram.memory[102][4] ),
    .I3(\u_cpu.rf_ram.memory[103][4] ),
    .S0(_01934_),
    .S1(_01648_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06505_ (.A1(_01646_),
    .A2(_02149_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06506_ (.I0(\u_cpu.rf_ram.memory[96][4] ),
    .I1(\u_cpu.rf_ram.memory[97][4] ),
    .I2(\u_cpu.rf_ram.memory[98][4] ),
    .I3(\u_cpu.rf_ram.memory[99][4] ),
    .S0(_01938_),
    .S1(_01824_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06507_ (.A1(_01937_),
    .A2(_02151_),
    .B(_01596_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06508_ (.I0(\u_cpu.rf_ram.memory[108][4] ),
    .I1(\u_cpu.rf_ram.memory[109][4] ),
    .I2(\u_cpu.rf_ram.memory[110][4] ),
    .I3(\u_cpu.rf_ram.memory[111][4] ),
    .S0(_02052_),
    .S1(_01827_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06509_ (.A1(_01941_),
    .A2(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06510_ (.I0(\u_cpu.rf_ram.memory[104][4] ),
    .I1(\u_cpu.rf_ram.memory[105][4] ),
    .I2(\u_cpu.rf_ram.memory[106][4] ),
    .I3(\u_cpu.rf_ram.memory[107][4] ),
    .S0(_02056_),
    .S1(_01624_),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06511_ (.A1(_02055_),
    .A2(_02155_),
    .B(_02058_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06512_ (.A1(_02150_),
    .A2(_02152_),
    .B1(_02154_),
    .B2(_02156_),
    .C(_01832_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06513_ (.I0(\u_cpu.rf_ram.memory[124][4] ),
    .I1(\u_cpu.rf_ram.memory[125][4] ),
    .I2(\u_cpu.rf_ram.memory[126][4] ),
    .I3(\u_cpu.rf_ram.memory[127][4] ),
    .S0(_01947_),
    .S1(_01669_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06514_ (.A1(_01582_),
    .A2(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06515_ (.I0(\u_cpu.rf_ram.memory[120][4] ),
    .I1(\u_cpu.rf_ram.memory[121][4] ),
    .I2(\u_cpu.rf_ram.memory[122][4] ),
    .I3(\u_cpu.rf_ram.memory[123][4] ),
    .S0(_01606_),
    .S1(_01837_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06516_ (.A1(_01836_),
    .A2(_02160_),
    .B(_01611_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06517_ (.I0(\u_cpu.rf_ram.memory[112][4] ),
    .I1(\u_cpu.rf_ram.memory[113][4] ),
    .I2(\u_cpu.rf_ram.memory[114][4] ),
    .I3(\u_cpu.rf_ram.memory[115][4] ),
    .S0(_02066_),
    .S1(_01840_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06518_ (.A1(_02065_),
    .A2(_02162_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06519_ (.I0(\u_cpu.rf_ram.memory[116][4] ),
    .I1(\u_cpu.rf_ram.memory[117][4] ),
    .I2(\u_cpu.rf_ram.memory[118][4] ),
    .I3(\u_cpu.rf_ram.memory[119][4] ),
    .S0(_02069_),
    .S1(_01685_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06520_ (.A1(_01683_),
    .A2(_02164_),
    .B(_01687_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06521_ (.A1(_02159_),
    .A2(_02161_),
    .B1(_02163_),
    .B2(_02165_),
    .C(_02072_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06522_ (.A1(_01580_),
    .A2(_02157_),
    .A3(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06523_ (.I0(\u_cpu.rf_ram.memory[92][4] ),
    .I1(\u_cpu.rf_ram.memory[93][4] ),
    .I2(\u_cpu.rf_ram.memory[94][4] ),
    .I3(\u_cpu.rf_ram.memory[95][4] ),
    .S0(_02075_),
    .S1(_01847_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06524_ (.A1(_01693_),
    .A2(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06525_ (.I0(\u_cpu.rf_ram.memory[88][4] ),
    .I1(\u_cpu.rf_ram.memory[89][4] ),
    .I2(\u_cpu.rf_ram.memory[90][4] ),
    .I3(\u_cpu.rf_ram.memory[91][4] ),
    .S0(_01961_),
    .S1(_01674_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06526_ (.A1(_01672_),
    .A2(_02170_),
    .B(_01963_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06527_ (.I0(\u_cpu.rf_ram.memory[80][4] ),
    .I1(\u_cpu.rf_ram.memory[81][4] ),
    .I2(\u_cpu.rf_ram.memory[82][4] ),
    .I3(\u_cpu.rf_ram.memory[83][4] ),
    .S0(_01584_),
    .S1(_01965_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06528_ (.A1(_01852_),
    .A2(_02172_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06529_ (.I0(\u_cpu.rf_ram.memory[84][4] ),
    .I1(\u_cpu.rf_ram.memory[85][4] ),
    .I2(\u_cpu.rf_ram.memory[86][4] ),
    .I3(\u_cpu.rf_ram.memory[87][4] ),
    .S0(_01855_),
    .S1(_02083_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06530_ (.A1(_02082_),
    .A2(_02174_),
    .B(_02085_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06531_ (.A1(_02169_),
    .A2(_02171_),
    .B1(_02173_),
    .B2(_02175_),
    .C(_01858_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06532_ (.I0(\u_cpu.rf_ram.memory[64][4] ),
    .I1(\u_cpu.rf_ram.memory[65][4] ),
    .I2(\u_cpu.rf_ram.memory[66][4] ),
    .I3(\u_cpu.rf_ram.memory[67][4] ),
    .S0(_01731_),
    .S1(_01972_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06533_ (.A1(_01971_),
    .A2(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06534_ (.I0(\u_cpu.rf_ram.memory[68][4] ),
    .I1(\u_cpu.rf_ram.memory[69][4] ),
    .I2(\u_cpu.rf_ram.memory[70][4] ),
    .I3(\u_cpu.rf_ram.memory[71][4] ),
    .S0(_01712_),
    .S1(_01863_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06535_ (.A1(_01862_),
    .A2(_02179_),
    .B(_01865_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06536_ (.I0(\u_cpu.rf_ram.memory[72][4] ),
    .I1(\u_cpu.rf_ram.memory[73][4] ),
    .I2(\u_cpu.rf_ram.memory[74][4] ),
    .I3(\u_cpu.rf_ram.memory[75][4] ),
    .S0(_01867_),
    .S1(_01695_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06537_ (.A1(_01705_),
    .A2(_02181_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06538_ (.I0(\u_cpu.rf_ram.memory[76][4] ),
    .I1(\u_cpu.rf_ram.memory[77][4] ),
    .I2(\u_cpu.rf_ram.memory[78][4] ),
    .I3(\u_cpu.rf_ram.memory[79][4] ),
    .S0(_01979_),
    .S1(_01726_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06539_ (.A1(_01724_),
    .A2(_02183_),
    .B(_01738_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06540_ (.A1(_02178_),
    .A2(_02180_),
    .B1(_02182_),
    .B2(_02184_),
    .C(_01982_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06541_ (.A1(_01958_),
    .A2(_02176_),
    .A3(_02185_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06542_ (.A1(_02167_),
    .A2(_02186_),
    .B(_01743_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06543_ (.I(_01538_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06544_ (.I0(\u_cpu.rf_ram.memory[136][4] ),
    .I1(\u_cpu.rf_ram.memory[137][4] ),
    .I2(\u_cpu.rf_ram.memory[138][4] ),
    .I3(\u_cpu.rf_ram.memory[139][4] ),
    .S0(_01747_),
    .S1(_01875_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06545_ (.A1(_02188_),
    .A2(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06546_ (.I0(\u_cpu.rf_ram.memory[140][4] ),
    .I1(\u_cpu.rf_ram.memory[141][4] ),
    .I2(\u_cpu.rf_ram.memory[142][4] ),
    .I3(\u_cpu.rf_ram.memory[143][4] ),
    .S0(_02101_),
    .S1(_01749_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06547_ (.A1(_01752_),
    .A2(_02191_),
    .B(_01756_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06548_ (.I0(\u_cpu.rf_ram.memory[128][4] ),
    .I1(\u_cpu.rf_ram.memory[129][4] ),
    .I2(\u_cpu.rf_ram.memory[130][4] ),
    .I3(\u_cpu.rf_ram.memory[131][4] ),
    .S0(_01542_),
    .S1(_01760_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06549_ (.A1(_01758_),
    .A2(_02193_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06550_ (.I0(\u_cpu.rf_ram.memory[132][4] ),
    .I1(\u_cpu.rf_ram.memory[133][4] ),
    .I2(\u_cpu.rf_ram.memory[134][4] ),
    .I3(\u_cpu.rf_ram.memory[135][4] ),
    .S0(_01993_),
    .S1(_02106_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06551_ (.A1(_01992_),
    .A2(_02195_),
    .B(_01574_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06552_ (.A1(_02190_),
    .A2(_02192_),
    .B1(_02194_),
    .B2(_02196_),
    .C(_01768_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06553_ (.A1(_02187_),
    .A2(_02197_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06554_ (.A1(_01497_),
    .A2(_02148_),
    .B(_02198_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06555_ (.I0(\u_cpu.rf_ram.memory[28][5] ),
    .I1(\u_cpu.rf_ram.memory[29][5] ),
    .I2(\u_cpu.rf_ram.memory[30][5] ),
    .I3(\u_cpu.rf_ram.memory[31][5] ),
    .S0(_01524_),
    .S1(_01771_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06556_ (.A1(_01523_),
    .A2(_02199_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06557_ (.I0(\u_cpu.rf_ram.memory[24][5] ),
    .I1(\u_cpu.rf_ram.memory[25][5] ),
    .I2(\u_cpu.rf_ram.memory[26][5] ),
    .I3(\u_cpu.rf_ram.memory[27][5] ),
    .S0(_01746_),
    .S1(_01774_),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06558_ (.A1(_01719_),
    .A2(_02201_),
    .B(_02001_),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06559_ (.I0(\u_cpu.rf_ram.memory[20][5] ),
    .I1(\u_cpu.rf_ram.memory[21][5] ),
    .I2(\u_cpu.rf_ram.memory[22][5] ),
    .I3(\u_cpu.rf_ram.memory[23][5] ),
    .S0(_01891_),
    .S1(_02003_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06560_ (.A1(_01890_),
    .A2(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06561_ (.I0(\u_cpu.rf_ram.memory[16][5] ),
    .I1(\u_cpu.rf_ram.memory[17][5] ),
    .I2(\u_cpu.rf_ram.memory[18][5] ),
    .I3(\u_cpu.rf_ram.memory[19][5] ),
    .S0(_02007_),
    .S1(_01518_),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06562_ (.A1(_02006_),
    .A2(_02205_),
    .B(_01728_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06563_ (.A1(_02200_),
    .A2(_02202_),
    .B1(_02204_),
    .B2(_02206_),
    .C(_01717_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06564_ (.I0(\u_cpu.rf_ram.memory[4][5] ),
    .I1(\u_cpu.rf_ram.memory[5][5] ),
    .I2(\u_cpu.rf_ram.memory[6][5] ),
    .I3(\u_cpu.rf_ram.memory[7][5] ),
    .S0(_01782_),
    .S1(_01897_),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06565_ (.A1(_02011_),
    .A2(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06566_ (.I0(\u_cpu.rf_ram.memory[0][5] ),
    .I1(\u_cpu.rf_ram.memory[1][5] ),
    .I2(\u_cpu.rf_ram.memory[2][5] ),
    .I3(\u_cpu.rf_ram.memory[3][5] ),
    .S0(_01786_),
    .S1(_01900_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06567_ (.A1(_01785_),
    .A2(_02210_),
    .B(_01902_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06568_ (.I0(\u_cpu.rf_ram.memory[8][5] ),
    .I1(\u_cpu.rf_ram.memory[9][5] ),
    .I2(\u_cpu.rf_ram.memory[10][5] ),
    .I3(\u_cpu.rf_ram.memory[11][5] ),
    .S0(_02016_),
    .S1(_01507_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06569_ (.A1(_01547_),
    .A2(_02212_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06570_ (.I0(\u_cpu.rf_ram.memory[12][5] ),
    .I1(\u_cpu.rf_ram.memory[13][5] ),
    .I2(\u_cpu.rf_ram.memory[14][5] ),
    .I3(\u_cpu.rf_ram.memory[15][5] ),
    .S0(_01550_),
    .S1(_01553_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06571_ (.A1(_01468_),
    .A2(_02214_),
    .B(_01792_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06572_ (.A1(_02209_),
    .A2(_02211_),
    .B1(_02213_),
    .B2(_02215_),
    .C(_01740_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06573_ (.I0(\u_cpu.rf_ram.memory[36][5] ),
    .I1(\u_cpu.rf_ram.memory[37][5] ),
    .I2(\u_cpu.rf_ram.memory[38][5] ),
    .I3(\u_cpu.rf_ram.memory[39][5] ),
    .S0(_01797_),
    .S1(_01680_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06574_ (.A1(_01796_),
    .A2(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06575_ (.I0(\u_cpu.rf_ram.memory[32][5] ),
    .I1(\u_cpu.rf_ram.memory[33][5] ),
    .I2(\u_cpu.rf_ram.memory[34][5] ),
    .I3(\u_cpu.rf_ram.memory[35][5] ),
    .S0(_01745_),
    .S1(_02024_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06576_ (.A1(_01559_),
    .A2(_02219_),
    .B(_01801_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06577_ (.I0(\u_cpu.rf_ram.memory[40][5] ),
    .I1(\u_cpu.rf_ram.memory[41][5] ),
    .I2(\u_cpu.rf_ram.memory[42][5] ),
    .I3(\u_cpu.rf_ram.memory[43][5] ),
    .S0(_02027_),
    .S1(_01563_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06578_ (.A1(_01634_),
    .A2(_02221_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06579_ (.I0(\u_cpu.rf_ram.memory[44][5] ),
    .I1(\u_cpu.rf_ram.memory[45][5] ),
    .I2(\u_cpu.rf_ram.memory[46][5] ),
    .I3(\u_cpu.rf_ram.memory[47][5] ),
    .S0(_01805_),
    .S1(_02030_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06580_ (.A1(_01915_),
    .A2(_02223_),
    .B(_01807_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06581_ (.A1(_02218_),
    .A2(_02220_),
    .B1(_02222_),
    .B2(_02224_),
    .C(_01665_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06582_ (.I0(\u_cpu.rf_ram.memory[60][5] ),
    .I1(\u_cpu.rf_ram.memory[61][5] ),
    .I2(\u_cpu.rf_ram.memory[62][5] ),
    .I3(\u_cpu.rf_ram.memory[63][5] ),
    .S0(_01668_),
    .S1(_02034_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06583_ (.A1(_01919_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06584_ (.I0(\u_cpu.rf_ram.memory[56][5] ),
    .I1(\u_cpu.rf_ram.memory[57][5] ),
    .I2(\u_cpu.rf_ram.memory[58][5] ),
    .I3(\u_cpu.rf_ram.memory[59][5] ),
    .S0(_01652_),
    .S1(_01812_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06585_ (.A1(_01651_),
    .A2(_02228_),
    .B(_01520_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06586_ (.I0(\u_cpu.rf_ram.memory[52][5] ),
    .I1(\u_cpu.rf_ram.memory[53][5] ),
    .I2(\u_cpu.rf_ram.memory[54][5] ),
    .I3(\u_cpu.rf_ram.memory[55][5] ),
    .S0(_01647_),
    .S1(_02040_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06587_ (.A1(_02039_),
    .A2(_02230_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06588_ (.I0(\u_cpu.rf_ram.memory[48][5] ),
    .I1(\u_cpu.rf_ram.memory[49][5] ),
    .I2(\u_cpu.rf_ram.memory[50][5] ),
    .I3(\u_cpu.rf_ram.memory[51][5] ),
    .S0(_01699_),
    .S1(_01927_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06589_ (.A1(_01926_),
    .A2(_02232_),
    .B(_01929_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06590_ (.A1(_02227_),
    .A2(_02229_),
    .B1(_02231_),
    .B2(_02233_),
    .C(_01489_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06591_ (.A1(_01795_),
    .A2(_02225_),
    .A3(_02234_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06592_ (.A1(_01692_),
    .A2(_02207_),
    .A3(_02216_),
    .B(_02235_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06593_ (.I0(\u_cpu.rf_ram.memory[100][5] ),
    .I1(\u_cpu.rf_ram.memory[101][5] ),
    .I2(\u_cpu.rf_ram.memory[102][5] ),
    .I3(\u_cpu.rf_ram.memory[103][5] ),
    .S0(_01934_),
    .S1(_01543_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06594_ (.A1(_01656_),
    .A2(_02237_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06595_ (.I0(\u_cpu.rf_ram.memory[96][5] ),
    .I1(\u_cpu.rf_ram.memory[97][5] ),
    .I2(\u_cpu.rf_ram.memory[98][5] ),
    .I3(\u_cpu.rf_ram.memory[99][5] ),
    .S0(_01938_),
    .S1(_01824_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06596_ (.A1(_01937_),
    .A2(_02239_),
    .B(_01596_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06597_ (.I0(\u_cpu.rf_ram.memory[108][5] ),
    .I1(\u_cpu.rf_ram.memory[109][5] ),
    .I2(\u_cpu.rf_ram.memory[110][5] ),
    .I3(\u_cpu.rf_ram.memory[111][5] ),
    .S0(_02052_),
    .S1(_01827_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06598_ (.A1(_01941_),
    .A2(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06599_ (.I0(\u_cpu.rf_ram.memory[104][5] ),
    .I1(\u_cpu.rf_ram.memory[105][5] ),
    .I2(\u_cpu.rf_ram.memory[106][5] ),
    .I3(\u_cpu.rf_ram.memory[107][5] ),
    .S0(_02056_),
    .S1(_01624_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06600_ (.A1(_02055_),
    .A2(_02243_),
    .B(_02058_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06601_ (.A1(_02238_),
    .A2(_02240_),
    .B1(_02242_),
    .B2(_02244_),
    .C(_01832_),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06602_ (.I0(\u_cpu.rf_ram.memory[124][5] ),
    .I1(\u_cpu.rf_ram.memory[125][5] ),
    .I2(\u_cpu.rf_ram.memory[126][5] ),
    .I3(\u_cpu.rf_ram.memory[127][5] ),
    .S0(_01947_),
    .S1(_01707_),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06603_ (.A1(_01582_),
    .A2(_02246_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06604_ (.I0(\u_cpu.rf_ram.memory[120][5] ),
    .I1(\u_cpu.rf_ram.memory[121][5] ),
    .I2(\u_cpu.rf_ram.memory[122][5] ),
    .I3(\u_cpu.rf_ram.memory[123][5] ),
    .S0(_01606_),
    .S1(_01837_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06605_ (.A1(_01836_),
    .A2(_02248_),
    .B(_01611_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06606_ (.I0(\u_cpu.rf_ram.memory[112][5] ),
    .I1(\u_cpu.rf_ram.memory[113][5] ),
    .I2(\u_cpu.rf_ram.memory[114][5] ),
    .I3(\u_cpu.rf_ram.memory[115][5] ),
    .S0(_02066_),
    .S1(_01840_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06607_ (.A1(_02065_),
    .A2(_02250_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06608_ (.I0(\u_cpu.rf_ram.memory[116][5] ),
    .I1(\u_cpu.rf_ram.memory[117][5] ),
    .I2(\u_cpu.rf_ram.memory[118][5] ),
    .I3(\u_cpu.rf_ram.memory[119][5] ),
    .S0(_02069_),
    .S1(_01638_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06609_ (.A1(_01604_),
    .A2(_02252_),
    .B(_01640_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06610_ (.A1(_02247_),
    .A2(_02249_),
    .B1(_02251_),
    .B2(_02253_),
    .C(_02072_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06611_ (.A1(_01580_),
    .A2(_02245_),
    .A3(_02254_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06612_ (.I0(\u_cpu.rf_ram.memory[92][5] ),
    .I1(\u_cpu.rf_ram.memory[93][5] ),
    .I2(\u_cpu.rf_ram.memory[94][5] ),
    .I3(\u_cpu.rf_ram.memory[95][5] ),
    .S0(_02075_),
    .S1(_01847_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06613_ (.A1(_01615_),
    .A2(_02256_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06614_ (.I0(\u_cpu.rf_ram.memory[88][5] ),
    .I1(\u_cpu.rf_ram.memory[89][5] ),
    .I2(\u_cpu.rf_ram.memory[90][5] ),
    .I3(\u_cpu.rf_ram.memory[91][5] ),
    .S0(_01961_),
    .S1(_01674_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06615_ (.A1(_01672_),
    .A2(_02258_),
    .B(_01963_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06616_ (.I0(\u_cpu.rf_ram.memory[80][5] ),
    .I1(\u_cpu.rf_ram.memory[81][5] ),
    .I2(\u_cpu.rf_ram.memory[82][5] ),
    .I3(\u_cpu.rf_ram.memory[83][5] ),
    .S0(_01584_),
    .S1(_01965_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06617_ (.A1(_01852_),
    .A2(_02260_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06618_ (.I0(\u_cpu.rf_ram.memory[84][5] ),
    .I1(\u_cpu.rf_ram.memory[85][5] ),
    .I2(\u_cpu.rf_ram.memory[86][5] ),
    .I3(\u_cpu.rf_ram.memory[87][5] ),
    .S0(_01855_),
    .S1(_02083_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06619_ (.A1(_02082_),
    .A2(_02262_),
    .B(_02085_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06620_ (.A1(_02257_),
    .A2(_02259_),
    .B1(_02261_),
    .B2(_02263_),
    .C(_01858_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06621_ (.I0(\u_cpu.rf_ram.memory[64][5] ),
    .I1(\u_cpu.rf_ram.memory[65][5] ),
    .I2(\u_cpu.rf_ram.memory[66][5] ),
    .I3(\u_cpu.rf_ram.memory[67][5] ),
    .S0(_01731_),
    .S1(_01972_),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06622_ (.A1(_01971_),
    .A2(_02265_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06623_ (.I0(\u_cpu.rf_ram.memory[68][5] ),
    .I1(\u_cpu.rf_ram.memory[69][5] ),
    .I2(\u_cpu.rf_ram.memory[70][5] ),
    .I3(\u_cpu.rf_ram.memory[71][5] ),
    .S0(_01712_),
    .S1(_01863_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06624_ (.A1(_01862_),
    .A2(_02267_),
    .B(_01865_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06625_ (.I0(\u_cpu.rf_ram.memory[72][5] ),
    .I1(\u_cpu.rf_ram.memory[73][5] ),
    .I2(\u_cpu.rf_ram.memory[74][5] ),
    .I3(\u_cpu.rf_ram.memory[75][5] ),
    .S0(_01867_),
    .S1(_01695_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06626_ (.A1(_01705_),
    .A2(_02269_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06627_ (.I0(\u_cpu.rf_ram.memory[76][5] ),
    .I1(\u_cpu.rf_ram.memory[77][5] ),
    .I2(\u_cpu.rf_ram.memory[78][5] ),
    .I3(\u_cpu.rf_ram.memory[79][5] ),
    .S0(_01979_),
    .S1(_01726_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06628_ (.A1(_01724_),
    .A2(_02271_),
    .B(_01702_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06629_ (.A1(_02266_),
    .A2(_02268_),
    .B1(_02270_),
    .B2(_02272_),
    .C(_01982_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06630_ (.A1(_01958_),
    .A2(_02264_),
    .A3(_02273_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06631_ (.A1(_02255_),
    .A2(_02274_),
    .B(_01475_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06632_ (.I0(\u_cpu.rf_ram.memory[136][5] ),
    .I1(\u_cpu.rf_ram.memory[137][5] ),
    .I2(\u_cpu.rf_ram.memory[138][5] ),
    .I3(\u_cpu.rf_ram.memory[139][5] ),
    .S0(_01764_),
    .S1(_01875_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06633_ (.A1(_02188_),
    .A2(_02276_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06634_ (.I0(\u_cpu.rf_ram.memory[140][5] ),
    .I1(\u_cpu.rf_ram.memory[141][5] ),
    .I2(\u_cpu.rf_ram.memory[142][5] ),
    .I3(\u_cpu.rf_ram.memory[143][5] ),
    .S0(_02101_),
    .S1(_01749_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06635_ (.A1(_01763_),
    .A2(_02278_),
    .B(_01756_),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06636_ (.I0(\u_cpu.rf_ram.memory[128][5] ),
    .I1(\u_cpu.rf_ram.memory[129][5] ),
    .I2(\u_cpu.rf_ram.memory[130][5] ),
    .I3(\u_cpu.rf_ram.memory[131][5] ),
    .S0(_01542_),
    .S1(_01544_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06637_ (.A1(_01539_),
    .A2(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06638_ (.I0(\u_cpu.rf_ram.memory[132][5] ),
    .I1(\u_cpu.rf_ram.memory[133][5] ),
    .I2(\u_cpu.rf_ram.memory[134][5] ),
    .I3(\u_cpu.rf_ram.memory[135][5] ),
    .S0(_01993_),
    .S1(_02106_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06639_ (.A1(_01992_),
    .A2(_02282_),
    .B(_01574_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06640_ (.A1(_02277_),
    .A2(_02279_),
    .B1(_02281_),
    .B2(_02283_),
    .C(_01470_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06641_ (.A1(_02275_),
    .A2(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06642_ (.A1(_01476_),
    .A2(_02236_),
    .B(_02285_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06643_ (.I0(\u_cpu.rf_ram.memory[28][6] ),
    .I1(\u_cpu.rf_ram.memory[29][6] ),
    .I2(\u_cpu.rf_ram.memory[30][6] ),
    .I3(\u_cpu.rf_ram.memory[31][6] ),
    .S0(_01524_),
    .S1(_01525_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06644_ (.A1(_01523_),
    .A2(_02286_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06645_ (.I0(\u_cpu.rf_ram.memory[24][6] ),
    .I1(\u_cpu.rf_ram.memory[25][6] ),
    .I2(\u_cpu.rf_ram.memory[26][6] ),
    .I3(\u_cpu.rf_ram.memory[27][6] ),
    .S0(_01746_),
    .S1(_01748_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06646_ (.A1(_01719_),
    .A2(_02288_),
    .B(_02001_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06647_ (.I0(\u_cpu.rf_ram.memory[20][6] ),
    .I1(\u_cpu.rf_ram.memory[21][6] ),
    .I2(\u_cpu.rf_ram.memory[22][6] ),
    .I3(\u_cpu.rf_ram.memory[23][6] ),
    .S0(_01891_),
    .S1(_02003_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06648_ (.A1(_01890_),
    .A2(_02290_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06649_ (.I0(\u_cpu.rf_ram.memory[16][6] ),
    .I1(\u_cpu.rf_ram.memory[17][6] ),
    .I2(\u_cpu.rf_ram.memory[18][6] ),
    .I3(\u_cpu.rf_ram.memory[19][6] ),
    .S0(_02007_),
    .S1(_01518_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06650_ (.A1(_02006_),
    .A2(_02292_),
    .B(_01728_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06651_ (.A1(_02287_),
    .A2(_02289_),
    .B1(_02291_),
    .B2(_02293_),
    .C(_01717_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06652_ (.I0(\u_cpu.rf_ram.memory[4][6] ),
    .I1(\u_cpu.rf_ram.memory[5][6] ),
    .I2(\u_cpu.rf_ram.memory[6][6] ),
    .I3(\u_cpu.rf_ram.memory[7][6] ),
    .S0(_01561_),
    .S1(_01897_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06653_ (.A1(_02011_),
    .A2(_02295_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06654_ (.I0(\u_cpu.rf_ram.memory[0][6] ),
    .I1(\u_cpu.rf_ram.memory[1][6] ),
    .I2(\u_cpu.rf_ram.memory[2][6] ),
    .I3(\u_cpu.rf_ram.memory[3][6] ),
    .S0(_01529_),
    .S1(_01900_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06655_ (.A1(_01528_),
    .A2(_02297_),
    .B(_01902_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06656_ (.I0(\u_cpu.rf_ram.memory[8][6] ),
    .I1(\u_cpu.rf_ram.memory[9][6] ),
    .I2(\u_cpu.rf_ram.memory[10][6] ),
    .I3(\u_cpu.rf_ram.memory[11][6] ),
    .S0(_02016_),
    .S1(_01507_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06657_ (.A1(_01547_),
    .A2(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06658_ (.I0(\u_cpu.rf_ram.memory[12][6] ),
    .I1(\u_cpu.rf_ram.memory[13][6] ),
    .I2(\u_cpu.rf_ram.memory[14][6] ),
    .I3(\u_cpu.rf_ram.memory[15][6] ),
    .S0(_01550_),
    .S1(_01553_),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06659_ (.A1(_01468_),
    .A2(_02301_),
    .B(_01521_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06660_ (.A1(_02296_),
    .A2(_02298_),
    .B1(_02300_),
    .B2(_02302_),
    .C(_01740_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06661_ (.I0(\u_cpu.rf_ram.memory[36][6] ),
    .I1(\u_cpu.rf_ram.memory[37][6] ),
    .I2(\u_cpu.rf_ram.memory[38][6] ),
    .I3(\u_cpu.rf_ram.memory[39][6] ),
    .S0(_01679_),
    .S1(_01680_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06662_ (.A1(_01629_),
    .A2(_02304_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06663_ (.I0(\u_cpu.rf_ram.memory[32][6] ),
    .I1(\u_cpu.rf_ram.memory[33][6] ),
    .I2(\u_cpu.rf_ram.memory[34][6] ),
    .I3(\u_cpu.rf_ram.memory[35][6] ),
    .S0(_01745_),
    .S1(_02024_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06664_ (.A1(_01559_),
    .A2(_02306_),
    .B(_01533_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06665_ (.I0(\u_cpu.rf_ram.memory[40][6] ),
    .I1(\u_cpu.rf_ram.memory[41][6] ),
    .I2(\u_cpu.rf_ram.memory[42][6] ),
    .I3(\u_cpu.rf_ram.memory[43][6] ),
    .S0(_02027_),
    .S1(_01563_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06666_ (.A1(_01634_),
    .A2(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06667_ (.I0(\u_cpu.rf_ram.memory[44][6] ),
    .I1(\u_cpu.rf_ram.memory[45][6] ),
    .I2(\u_cpu.rf_ram.memory[46][6] ),
    .I3(\u_cpu.rf_ram.memory[47][6] ),
    .S0(_01661_),
    .S1(_02030_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06668_ (.A1(_01915_),
    .A2(_02310_),
    .B(_01663_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06669_ (.A1(_02305_),
    .A2(_02307_),
    .B1(_02309_),
    .B2(_02311_),
    .C(_01665_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06670_ (.I0(\u_cpu.rf_ram.memory[60][6] ),
    .I1(\u_cpu.rf_ram.memory[61][6] ),
    .I2(\u_cpu.rf_ram.memory[62][6] ),
    .I3(\u_cpu.rf_ram.memory[63][6] ),
    .S0(_01668_),
    .S1(_02034_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06671_ (.A1(_01919_),
    .A2(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06672_ (.I0(\u_cpu.rf_ram.memory[56][6] ),
    .I1(\u_cpu.rf_ram.memory[57][6] ),
    .I2(\u_cpu.rf_ram.memory[58][6] ),
    .I3(\u_cpu.rf_ram.memory[59][6] ),
    .S0(_01652_),
    .S1(_01552_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06673_ (.A1(_01651_),
    .A2(_02315_),
    .B(_01520_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06674_ (.I0(\u_cpu.rf_ram.memory[52][6] ),
    .I1(\u_cpu.rf_ram.memory[53][6] ),
    .I2(\u_cpu.rf_ram.memory[54][6] ),
    .I3(\u_cpu.rf_ram.memory[55][6] ),
    .S0(_01647_),
    .S1(_02040_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06675_ (.A1(_02039_),
    .A2(_02317_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06676_ (.I0(\u_cpu.rf_ram.memory[48][6] ),
    .I1(\u_cpu.rf_ram.memory[49][6] ),
    .I2(\u_cpu.rf_ram.memory[50][6] ),
    .I3(\u_cpu.rf_ram.memory[51][6] ),
    .S0(_01699_),
    .S1(_01927_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06677_ (.A1(_01926_),
    .A2(_02319_),
    .B(_01929_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06678_ (.A1(_02314_),
    .A2(_02316_),
    .B1(_02318_),
    .B2(_02320_),
    .C(_01489_),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06679_ (.A1(_01493_),
    .A2(_02312_),
    .A3(_02321_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06680_ (.A1(_01692_),
    .A2(_02294_),
    .A3(_02303_),
    .B(_02322_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06681_ (.I0(\u_cpu.rf_ram.memory[100][6] ),
    .I1(\u_cpu.rf_ram.memory[101][6] ),
    .I2(\u_cpu.rf_ram.memory[102][6] ),
    .I3(\u_cpu.rf_ram.memory[103][6] ),
    .S0(_01934_),
    .S1(_01543_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06682_ (.A1(_01656_),
    .A2(_02324_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06683_ (.I0(\u_cpu.rf_ram.memory[96][6] ),
    .I1(\u_cpu.rf_ram.memory[97][6] ),
    .I2(\u_cpu.rf_ram.memory[98][6] ),
    .I3(\u_cpu.rf_ram.memory[99][6] ),
    .S0(_01938_),
    .S1(_01593_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06684_ (.A1(_01937_),
    .A2(_02326_),
    .B(_01596_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06685_ (.I0(\u_cpu.rf_ram.memory[108][6] ),
    .I1(\u_cpu.rf_ram.memory[109][6] ),
    .I2(\u_cpu.rf_ram.memory[110][6] ),
    .I3(\u_cpu.rf_ram.memory[111][6] ),
    .S0(_02052_),
    .S1(_01506_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06686_ (.A1(_01941_),
    .A2(_02328_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06687_ (.I0(\u_cpu.rf_ram.memory[104][6] ),
    .I1(\u_cpu.rf_ram.memory[105][6] ),
    .I2(\u_cpu.rf_ram.memory[106][6] ),
    .I3(\u_cpu.rf_ram.memory[107][6] ),
    .S0(_02056_),
    .S1(_01624_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06688_ (.A1(_02055_),
    .A2(_02330_),
    .B(_02058_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06689_ (.A1(_02325_),
    .A2(_02327_),
    .B1(_02329_),
    .B2(_02331_),
    .C(_01577_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06690_ (.I0(\u_cpu.rf_ram.memory[124][6] ),
    .I1(\u_cpu.rf_ram.memory[125][6] ),
    .I2(\u_cpu.rf_ram.memory[126][6] ),
    .I3(\u_cpu.rf_ram.memory[127][6] ),
    .S0(_01947_),
    .S1(_01707_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06691_ (.A1(_01582_),
    .A2(_02333_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06692_ (.I0(\u_cpu.rf_ram.memory[120][6] ),
    .I1(\u_cpu.rf_ram.memory[121][6] ),
    .I2(\u_cpu.rf_ram.memory[122][6] ),
    .I3(\u_cpu.rf_ram.memory[123][6] ),
    .S0(_01606_),
    .S1(_01608_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06693_ (.A1(_01660_),
    .A2(_02335_),
    .B(_01611_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06694_ (.I0(\u_cpu.rf_ram.memory[112][6] ),
    .I1(\u_cpu.rf_ram.memory[113][6] ),
    .I2(\u_cpu.rf_ram.memory[114][6] ),
    .I3(\u_cpu.rf_ram.memory[115][6] ),
    .S0(_02066_),
    .S1(_01631_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06695_ (.A1(_02065_),
    .A2(_02337_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06696_ (.I0(\u_cpu.rf_ram.memory[116][6] ),
    .I1(\u_cpu.rf_ram.memory[117][6] ),
    .I2(\u_cpu.rf_ram.memory[118][6] ),
    .I3(\u_cpu.rf_ram.memory[119][6] ),
    .S0(_02069_),
    .S1(_01638_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06697_ (.A1(_01604_),
    .A2(_02339_),
    .B(_01640_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06698_ (.A1(_02334_),
    .A2(_02336_),
    .B1(_02338_),
    .B2(_02340_),
    .C(_02072_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06699_ (.A1(_01580_),
    .A2(_02332_),
    .A3(_02341_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06700_ (.I0(\u_cpu.rf_ram.memory[92][6] ),
    .I1(\u_cpu.rf_ram.memory[93][6] ),
    .I2(\u_cpu.rf_ram.memory[94][6] ),
    .I3(\u_cpu.rf_ram.memory[95][6] ),
    .S0(_02075_),
    .S1(_01619_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06701_ (.A1(_01615_),
    .A2(_02343_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06702_ (.I0(\u_cpu.rf_ram.memory[88][6] ),
    .I1(\u_cpu.rf_ram.memory[89][6] ),
    .I2(\u_cpu.rf_ram.memory[90][6] ),
    .I3(\u_cpu.rf_ram.memory[91][6] ),
    .S0(_01961_),
    .S1(_01674_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06703_ (.A1(_01672_),
    .A2(_02345_),
    .B(_01963_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06704_ (.I0(\u_cpu.rf_ram.memory[80][6] ),
    .I1(\u_cpu.rf_ram.memory[81][6] ),
    .I2(\u_cpu.rf_ram.memory[82][6] ),
    .I3(\u_cpu.rf_ram.memory[83][6] ),
    .S0(_01584_),
    .S1(_01965_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06705_ (.A1(_01678_),
    .A2(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06706_ (.I0(\u_cpu.rf_ram.memory[84][6] ),
    .I1(\u_cpu.rf_ram.memory[85][6] ),
    .I2(\u_cpu.rf_ram.memory[86][6] ),
    .I3(\u_cpu.rf_ram.memory[87][6] ),
    .S0(_01684_),
    .S1(_02083_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06707_ (.A1(_02082_),
    .A2(_02349_),
    .B(_02085_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06708_ (.A1(_02344_),
    .A2(_02346_),
    .B1(_02348_),
    .B2(_02350_),
    .C(_01689_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06709_ (.I0(\u_cpu.rf_ram.memory[64][6] ),
    .I1(\u_cpu.rf_ram.memory[65][6] ),
    .I2(\u_cpu.rf_ram.memory[66][6] ),
    .I3(\u_cpu.rf_ram.memory[67][6] ),
    .S0(_01731_),
    .S1(_01972_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06710_ (.A1(_01971_),
    .A2(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06711_ (.I0(\u_cpu.rf_ram.memory[68][6] ),
    .I1(\u_cpu.rf_ram.memory[69][6] ),
    .I2(\u_cpu.rf_ram.memory[70][6] ),
    .I3(\u_cpu.rf_ram.memory[71][6] ),
    .S0(_01712_),
    .S1(_01713_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06712_ (.A1(_01711_),
    .A2(_02354_),
    .B(_01715_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06713_ (.I0(\u_cpu.rf_ram.memory[72][6] ),
    .I1(\u_cpu.rf_ram.memory[73][6] ),
    .I2(\u_cpu.rf_ram.memory[74][6] ),
    .I3(\u_cpu.rf_ram.memory[75][6] ),
    .S0(_01694_),
    .S1(_01695_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06714_ (.A1(_01705_),
    .A2(_02356_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06715_ (.I0(\u_cpu.rf_ram.memory[76][6] ),
    .I1(\u_cpu.rf_ram.memory[77][6] ),
    .I2(\u_cpu.rf_ram.memory[78][6] ),
    .I3(\u_cpu.rf_ram.memory[79][6] ),
    .S0(_01979_),
    .S1(_01726_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06716_ (.A1(_01724_),
    .A2(_02358_),
    .B(_01702_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06717_ (.A1(_02353_),
    .A2(_02355_),
    .B1(_02357_),
    .B2(_02359_),
    .C(_01982_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06718_ (.A1(_01958_),
    .A2(_02351_),
    .A3(_02360_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06719_ (.A1(_02342_),
    .A2(_02361_),
    .B(_01475_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06720_ (.I0(\u_cpu.rf_ram.memory[128][6] ),
    .I1(\u_cpu.rf_ram.memory[129][6] ),
    .I2(\u_cpu.rf_ram.memory[130][6] ),
    .I3(\u_cpu.rf_ram.memory[131][6] ),
    .S0(_01764_),
    .S1(_01765_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06721_ (.A1(_02188_),
    .A2(_02363_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06722_ (.I0(\u_cpu.rf_ram.memory[132][6] ),
    .I1(\u_cpu.rf_ram.memory[133][6] ),
    .I2(\u_cpu.rf_ram.memory[134][6] ),
    .I3(\u_cpu.rf_ram.memory[135][6] ),
    .S0(_02101_),
    .S1(_01749_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06723_ (.A1(_01763_),
    .A2(_02365_),
    .B(_01485_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06724_ (.I0(\u_cpu.rf_ram.memory[136][6] ),
    .I1(\u_cpu.rf_ram.memory[137][6] ),
    .I2(\u_cpu.rf_ram.memory[138][6] ),
    .I3(\u_cpu.rf_ram.memory[139][6] ),
    .S0(_01542_),
    .S1(_01544_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06725_ (.A1(_01539_),
    .A2(_02367_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06726_ (.I0(\u_cpu.rf_ram.memory[140][6] ),
    .I1(\u_cpu.rf_ram.memory[141][6] ),
    .I2(\u_cpu.rf_ram.memory[142][6] ),
    .I3(\u_cpu.rf_ram.memory[143][6] ),
    .S0(_01993_),
    .S1(_02106_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06727_ (.A1(_01992_),
    .A2(_02369_),
    .B(_01556_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06728_ (.A1(_02364_),
    .A2(_02366_),
    .B1(_02368_),
    .B2(_02370_),
    .C(_01470_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06729_ (.A1(_02362_),
    .A2(_02371_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06730_ (.A1(_01476_),
    .A2(_02323_),
    .B(_02372_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06731_ (.I0(\u_cpu.rf_ram.memory[28][7] ),
    .I1(\u_cpu.rf_ram.memory[29][7] ),
    .I2(\u_cpu.rf_ram.memory[30][7] ),
    .I3(\u_cpu.rf_ram.memory[31][7] ),
    .S0(_01524_),
    .S1(_01525_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06732_ (.A1(_01523_),
    .A2(_02373_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06733_ (.I0(\u_cpu.rf_ram.memory[24][7] ),
    .I1(\u_cpu.rf_ram.memory[25][7] ),
    .I2(\u_cpu.rf_ram.memory[26][7] ),
    .I3(\u_cpu.rf_ram.memory[27][7] ),
    .S0(_01746_),
    .S1(_01748_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06734_ (.A1(_01719_),
    .A2(_02375_),
    .B(_02001_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06735_ (.I0(\u_cpu.rf_ram.memory[20][7] ),
    .I1(\u_cpu.rf_ram.memory[21][7] ),
    .I2(\u_cpu.rf_ram.memory[22][7] ),
    .I3(\u_cpu.rf_ram.memory[23][7] ),
    .S0(_01570_),
    .S1(_02003_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06736_ (.A1(_01567_),
    .A2(_02377_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06737_ (.I0(\u_cpu.rf_ram.memory[16][7] ),
    .I1(\u_cpu.rf_ram.memory[17][7] ),
    .I2(\u_cpu.rf_ram.memory[18][7] ),
    .I3(\u_cpu.rf_ram.memory[19][7] ),
    .S0(_02007_),
    .S1(_01518_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06738_ (.A1(_02006_),
    .A2(_02379_),
    .B(_01728_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06739_ (.A1(_02374_),
    .A2(_02376_),
    .B1(_02378_),
    .B2(_02380_),
    .C(_01717_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06740_ (.I0(\u_cpu.rf_ram.memory[4][7] ),
    .I1(\u_cpu.rf_ram.memory[5][7] ),
    .I2(\u_cpu.rf_ram.memory[6][7] ),
    .I3(\u_cpu.rf_ram.memory[7][7] ),
    .S0(_01561_),
    .S1(_01564_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06741_ (.A1(_02011_),
    .A2(_02382_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06742_ (.I0(\u_cpu.rf_ram.memory[0][7] ),
    .I1(\u_cpu.rf_ram.memory[1][7] ),
    .I2(\u_cpu.rf_ram.memory[2][7] ),
    .I3(\u_cpu.rf_ram.memory[3][7] ),
    .S0(_01529_),
    .S1(_01530_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06743_ (.A1(_01528_),
    .A2(_02384_),
    .B(_01534_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06744_ (.I0(\u_cpu.rf_ram.memory[8][7] ),
    .I1(\u_cpu.rf_ram.memory[9][7] ),
    .I2(\u_cpu.rf_ram.memory[10][7] ),
    .I3(\u_cpu.rf_ram.memory[11][7] ),
    .S0(_02016_),
    .S1(_01507_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06745_ (.A1(_01547_),
    .A2(_02386_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06746_ (.I0(\u_cpu.rf_ram.memory[12][7] ),
    .I1(\u_cpu.rf_ram.memory[13][7] ),
    .I2(\u_cpu.rf_ram.memory[14][7] ),
    .I3(\u_cpu.rf_ram.memory[15][7] ),
    .S0(_01550_),
    .S1(_01553_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06747_ (.A1(_01468_),
    .A2(_02388_),
    .B(_01521_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06748_ (.A1(_02383_),
    .A2(_02385_),
    .B1(_02387_),
    .B2(_02389_),
    .C(_01740_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06749_ (.I0(\u_cpu.rf_ram.memory[36][7] ),
    .I1(\u_cpu.rf_ram.memory[37][7] ),
    .I2(\u_cpu.rf_ram.memory[38][7] ),
    .I3(\u_cpu.rf_ram.memory[39][7] ),
    .S0(_01679_),
    .S1(_01680_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06750_ (.A1(_01629_),
    .A2(_02391_),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06751_ (.I0(\u_cpu.rf_ram.memory[32][7] ),
    .I1(\u_cpu.rf_ram.memory[33][7] ),
    .I2(\u_cpu.rf_ram.memory[34][7] ),
    .I3(\u_cpu.rf_ram.memory[35][7] ),
    .S0(_01745_),
    .S1(_02024_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06752_ (.A1(_01559_),
    .A2(_02393_),
    .B(_01533_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06753_ (.I0(\u_cpu.rf_ram.memory[40][7] ),
    .I1(\u_cpu.rf_ram.memory[41][7] ),
    .I2(\u_cpu.rf_ram.memory[42][7] ),
    .I3(\u_cpu.rf_ram.memory[43][7] ),
    .S0(_02027_),
    .S1(_01563_),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06754_ (.A1(_01634_),
    .A2(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06755_ (.I0(\u_cpu.rf_ram.memory[44][7] ),
    .I1(\u_cpu.rf_ram.memory[45][7] ),
    .I2(\u_cpu.rf_ram.memory[46][7] ),
    .I3(\u_cpu.rf_ram.memory[47][7] ),
    .S0(_01661_),
    .S1(_02030_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06756_ (.A1(_01538_),
    .A2(_02397_),
    .B(_01663_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06757_ (.A1(_02392_),
    .A2(_02394_),
    .B1(_02396_),
    .B2(_02398_),
    .C(_01665_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06758_ (.I0(\u_cpu.rf_ram.memory[60][7] ),
    .I1(\u_cpu.rf_ram.memory[61][7] ),
    .I2(\u_cpu.rf_ram.memory[62][7] ),
    .I3(\u_cpu.rf_ram.memory[63][7] ),
    .S0(_01668_),
    .S1(_02034_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06759_ (.A1(_01667_),
    .A2(_02400_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06760_ (.I0(\u_cpu.rf_ram.memory[56][7] ),
    .I1(\u_cpu.rf_ram.memory[57][7] ),
    .I2(\u_cpu.rf_ram.memory[58][7] ),
    .I3(\u_cpu.rf_ram.memory[59][7] ),
    .S0(_01652_),
    .S1(_01552_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06761_ (.A1(_01651_),
    .A2(_02402_),
    .B(_01520_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06762_ (.I0(\u_cpu.rf_ram.memory[52][7] ),
    .I1(\u_cpu.rf_ram.memory[53][7] ),
    .I2(\u_cpu.rf_ram.memory[54][7] ),
    .I3(\u_cpu.rf_ram.memory[55][7] ),
    .S0(_01647_),
    .S1(_02040_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06763_ (.A1(_02039_),
    .A2(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06764_ (.I0(\u_cpu.rf_ram.memory[48][7] ),
    .I1(\u_cpu.rf_ram.memory[49][7] ),
    .I2(\u_cpu.rf_ram.memory[50][7] ),
    .I3(\u_cpu.rf_ram.memory[51][7] ),
    .S0(_01699_),
    .S1(_01700_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06765_ (.A1(_01698_),
    .A2(_02406_),
    .B(_01654_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06766_ (.A1(_02401_),
    .A2(_02403_),
    .B1(_02405_),
    .B2(_02407_),
    .C(_01489_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06767_ (.A1(_01493_),
    .A2(_02399_),
    .A3(_02408_),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06768_ (.A1(_01692_),
    .A2(_02381_),
    .A3(_02390_),
    .B(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06769_ (.I0(\u_cpu.rf_ram.memory[100][7] ),
    .I1(\u_cpu.rf_ram.memory[101][7] ),
    .I2(\u_cpu.rf_ram.memory[102][7] ),
    .I3(\u_cpu.rf_ram.memory[103][7] ),
    .S0(_01569_),
    .S1(_01543_),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06770_ (.A1(_01656_),
    .A2(_02411_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06771_ (.I0(\u_cpu.rf_ram.memory[96][7] ),
    .I1(\u_cpu.rf_ram.memory[97][7] ),
    .I2(\u_cpu.rf_ram.memory[98][7] ),
    .I3(\u_cpu.rf_ram.memory[99][7] ),
    .S0(_01590_),
    .S1(_01593_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06772_ (.A1(_01589_),
    .A2(_02413_),
    .B(_01596_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06773_ (.I0(\u_cpu.rf_ram.memory[108][7] ),
    .I1(\u_cpu.rf_ram.memory[109][7] ),
    .I2(\u_cpu.rf_ram.memory[110][7] ),
    .I3(\u_cpu.rf_ram.memory[111][7] ),
    .S0(_02052_),
    .S1(_01506_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06774_ (.A1(_01735_),
    .A2(_02415_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06775_ (.I0(\u_cpu.rf_ram.memory[104][7] ),
    .I1(\u_cpu.rf_ram.memory[105][7] ),
    .I2(\u_cpu.rf_ram.memory[106][7] ),
    .I3(\u_cpu.rf_ram.memory[107][7] ),
    .S0(_02056_),
    .S1(_01624_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06776_ (.A1(_02055_),
    .A2(_02417_),
    .B(_02058_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06777_ (.A1(_02412_),
    .A2(_02414_),
    .B1(_02416_),
    .B2(_02418_),
    .C(_01577_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06778_ (.I0(\u_cpu.rf_ram.memory[124][7] ),
    .I1(\u_cpu.rf_ram.memory[125][7] ),
    .I2(\u_cpu.rf_ram.memory[126][7] ),
    .I3(\u_cpu.rf_ram.memory[127][7] ),
    .S0(_01706_),
    .S1(_01707_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06779_ (.A1(_01582_),
    .A2(_02420_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06780_ (.I0(\u_cpu.rf_ram.memory[120][7] ),
    .I1(\u_cpu.rf_ram.memory[121][7] ),
    .I2(\u_cpu.rf_ram.memory[122][7] ),
    .I3(\u_cpu.rf_ram.memory[123][7] ),
    .S0(_01606_),
    .S1(_01608_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06781_ (.A1(_01660_),
    .A2(_02422_),
    .B(_01611_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06782_ (.I0(\u_cpu.rf_ram.memory[112][7] ),
    .I1(\u_cpu.rf_ram.memory[113][7] ),
    .I2(\u_cpu.rf_ram.memory[114][7] ),
    .I3(\u_cpu.rf_ram.memory[115][7] ),
    .S0(_02066_),
    .S1(_01631_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06783_ (.A1(_02065_),
    .A2(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06784_ (.I0(\u_cpu.rf_ram.memory[116][7] ),
    .I1(\u_cpu.rf_ram.memory[117][7] ),
    .I2(\u_cpu.rf_ram.memory[118][7] ),
    .I3(\u_cpu.rf_ram.memory[119][7] ),
    .S0(_02069_),
    .S1(_01638_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06785_ (.A1(_01604_),
    .A2(_02426_),
    .B(_01640_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06786_ (.A1(_02421_),
    .A2(_02423_),
    .B1(_02425_),
    .B2(_02427_),
    .C(_02072_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06787_ (.A1(_01580_),
    .A2(_02419_),
    .A3(_02428_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06788_ (.I0(\u_cpu.rf_ram.memory[92][7] ),
    .I1(\u_cpu.rf_ram.memory[93][7] ),
    .I2(\u_cpu.rf_ram.memory[94][7] ),
    .I3(\u_cpu.rf_ram.memory[95][7] ),
    .S0(_02075_),
    .S1(_01619_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06789_ (.A1(_01615_),
    .A2(_02430_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06790_ (.I0(\u_cpu.rf_ram.memory[88][7] ),
    .I1(\u_cpu.rf_ram.memory[89][7] ),
    .I2(\u_cpu.rf_ram.memory[90][7] ),
    .I3(\u_cpu.rf_ram.memory[91][7] ),
    .S0(_01673_),
    .S1(_01674_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06791_ (.A1(_01672_),
    .A2(_02432_),
    .B(_01676_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06792_ (.I0(\u_cpu.rf_ram.memory[80][7] ),
    .I1(\u_cpu.rf_ram.memory[81][7] ),
    .I2(\u_cpu.rf_ram.memory[82][7] ),
    .I3(\u_cpu.rf_ram.memory[83][7] ),
    .S0(_01584_),
    .S1(_01586_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06793_ (.A1(_01678_),
    .A2(_02434_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06794_ (.I0(\u_cpu.rf_ram.memory[84][7] ),
    .I1(\u_cpu.rf_ram.memory[85][7] ),
    .I2(\u_cpu.rf_ram.memory[86][7] ),
    .I3(\u_cpu.rf_ram.memory[87][7] ),
    .S0(_01684_),
    .S1(_02083_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06795_ (.A1(_02082_),
    .A2(_02436_),
    .B(_02085_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06796_ (.A1(_02431_),
    .A2(_02433_),
    .B1(_02435_),
    .B2(_02437_),
    .C(_01689_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06797_ (.I0(\u_cpu.rf_ram.memory[64][7] ),
    .I1(\u_cpu.rf_ram.memory[65][7] ),
    .I2(\u_cpu.rf_ram.memory[66][7] ),
    .I3(\u_cpu.rf_ram.memory[67][7] ),
    .S0(_01731_),
    .S1(_01732_),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06798_ (.A1(_01730_),
    .A2(_02439_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06799_ (.I0(\u_cpu.rf_ram.memory[68][7] ),
    .I1(\u_cpu.rf_ram.memory[69][7] ),
    .I2(\u_cpu.rf_ram.memory[70][7] ),
    .I3(\u_cpu.rf_ram.memory[71][7] ),
    .S0(_01712_),
    .S1(_01713_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06800_ (.A1(_01711_),
    .A2(_02441_),
    .B(_01715_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06801_ (.I0(\u_cpu.rf_ram.memory[72][7] ),
    .I1(\u_cpu.rf_ram.memory[73][7] ),
    .I2(\u_cpu.rf_ram.memory[74][7] ),
    .I3(\u_cpu.rf_ram.memory[75][7] ),
    .S0(_01694_),
    .S1(_01695_),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06802_ (.A1(_01705_),
    .A2(_02443_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06803_ (.I0(\u_cpu.rf_ram.memory[76][7] ),
    .I1(\u_cpu.rf_ram.memory[77][7] ),
    .I2(\u_cpu.rf_ram.memory[78][7] ),
    .I3(\u_cpu.rf_ram.memory[79][7] ),
    .S0(_01725_),
    .S1(_01726_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06804_ (.A1(_01724_),
    .A2(_02445_),
    .B(_01702_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06805_ (.A1(_02440_),
    .A2(_02442_),
    .B1(_02444_),
    .B2(_02446_),
    .C(_01613_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06806_ (.A1(_01498_),
    .A2(_02438_),
    .A3(_02447_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06807_ (.A1(_02429_),
    .A2(_02448_),
    .B(_01475_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06808_ (.I0(\u_cpu.rf_ram.memory[128][7] ),
    .I1(\u_cpu.rf_ram.memory[129][7] ),
    .I2(\u_cpu.rf_ram.memory[130][7] ),
    .I3(\u_cpu.rf_ram.memory[131][7] ),
    .S0(_01764_),
    .S1(_01765_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06809_ (.A1(_02188_),
    .A2(_02450_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06810_ (.I0(\u_cpu.rf_ram.memory[132][7] ),
    .I1(\u_cpu.rf_ram.memory[133][7] ),
    .I2(\u_cpu.rf_ram.memory[134][7] ),
    .I3(\u_cpu.rf_ram.memory[135][7] ),
    .S0(_02101_),
    .S1(_01749_),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06811_ (.A1(_01763_),
    .A2(_02452_),
    .B(_01485_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06812_ (.I0(\u_cpu.rf_ram.memory[140][7] ),
    .I1(\u_cpu.rf_ram.memory[141][7] ),
    .I2(\u_cpu.rf_ram.memory[142][7] ),
    .I3(\u_cpu.rf_ram.memory[143][7] ),
    .S0(_01542_),
    .S1(_01544_),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06813_ (.A1(_01560_),
    .A2(_02454_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06814_ (.I0(\u_cpu.rf_ram.memory[136][7] ),
    .I1(\u_cpu.rf_ram.memory[137][7] ),
    .I2(\u_cpu.rf_ram.memory[138][7] ),
    .I3(\u_cpu.rf_ram.memory[139][7] ),
    .S0(_01759_),
    .S1(_02106_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06815_ (.A1(_02188_),
    .A2(_02456_),
    .B(_01556_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06816_ (.A1(_02451_),
    .A2(_02453_),
    .B1(_02455_),
    .B2(_02457_),
    .C(_01470_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06817_ (.A1(_02449_),
    .A2(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06818_ (.A1(_01476_),
    .A2(_02410_),
    .B(_02459_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06819_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06820_ (.I(_02460_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06821_ (.I(_02461_),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06822_ (.I(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06823_ (.A1(_01451_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06824_ (.A1(_02463_),
    .A2(\u_cpu.cpu.bufreg.i_sh_signed ),
    .B(_02464_),
    .C(_01444_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06825_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06826_ (.I(\u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06827_ (.A1(\u_cpu.cpu.decode.opcode[2] ),
    .A2(\u_cpu.cpu.decode.opcode[0] ),
    .A3(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06828_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_02467_),
    .A3(_02468_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06829_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_02468_),
    .B(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06830_ (.A1(_01443_),
    .A2(\u_cpu.cpu.branch_op ),
    .A3(\u_cpu.cpu.csr_d_sel ),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06831_ (.A1(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .A2(\u_cpu.cpu.immdec.imm31 ),
    .A3(_02471_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06832_ (.A1(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .A2(_02469_),
    .A3(_02470_),
    .B(_02472_),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06833_ (.I(\u_cpu.rf_ram.regzero ),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06834_ (.A1(\u_cpu.rf_ram.rdata[0] ),
    .A2(_02474_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06835_ (.A1(\u_cpu.rf_ram_if.rdata1[0] ),
    .A2(\u_cpu.rf_ram_if.rtrig1 ),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06836_ (.A1(\u_cpu.rf_ram_if.rtrig1 ),
    .A2(_02475_),
    .B(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06837_ (.I0(_02473_),
    .I1(_02477_),
    .S(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06838_ (.A1(_02465_),
    .A2(_02478_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06839_ (.I(\u_cpu.cpu.alu.i_rs1 ),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06840_ (.A1(_02480_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06841_ (.A1(_02466_),
    .A2(_02479_),
    .B(_02481_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06842_ (.A1(_02462_),
    .A2(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06843_ (.A1(_02462_),
    .A2(_02465_),
    .B(_02483_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06844_ (.I(_01463_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06845_ (.I(_01451_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06846_ (.A1(_02485_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06847_ (.I(_01452_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06848_ (.A1(_02487_),
    .A2(_01439_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06849_ (.A1(_02487_),
    .A2(_02480_),
    .B(_02488_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06850_ (.I(_01451_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06851_ (.I(_02490_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06852_ (.I(\u_cpu.cpu.bne_or_bge ),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06853_ (.I(_02492_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06854_ (.A1(_02491_),
    .A2(_02493_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06855_ (.I(_02485_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06856_ (.A1(_02495_),
    .A2(_02489_),
    .B(_02493_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06857_ (.A1(_01447_),
    .A2(_01450_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06858_ (.I(\u_cpu.cpu.state.o_cnt_r[3] ),
    .Z(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06859_ (.I(\u_cpu.cpu.decode.op22 ),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06860_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06861_ (.I(_02500_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06862_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_01447_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06863_ (.A1(_02498_),
    .A2(_02499_),
    .A3(_02501_),
    .A4(_02502_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06864_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06865_ (.I(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06866_ (.A1(_02505_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .B(_02500_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06867_ (.A1(_01448_),
    .A2(_01449_),
    .A3(_01446_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06868_ (.A1(_02460_),
    .A2(_02507_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06869_ (.A1(_02504_),
    .A2(_02501_),
    .B(_02506_),
    .C(_02508_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06870_ (.A1(_02497_),
    .A2(_02477_),
    .B1(_02503_),
    .B2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .C(_02509_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _06871_ (.A1(_02486_),
    .A2(_02489_),
    .A3(_02494_),
    .B1(_02496_),
    .B2(_02510_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06872_ (.A1(_02484_),
    .A2(_02511_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06873_ (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06874_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_01462_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06875_ (.I(_02514_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06876_ (.A1(_02513_),
    .A2(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06877_ (.A1(_02512_),
    .A2(_02516_),
    .ZN(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06878_ (.I(_01444_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06879_ (.I(_02517_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06880_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.init_done ),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06881_ (.A1(_02517_),
    .A2(_02514_),
    .A3(_02519_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06882_ (.I(\u_cpu.cpu.decode.opcode[0] ),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06883_ (.I(_01452_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06884_ (.A1(_02490_),
    .A2(_02522_),
    .B(_02464_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06885_ (.I(_01443_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06886_ (.A1(_02517_),
    .A2(_02521_),
    .A3(_02523_),
    .B(_02524_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06887_ (.A1(_02460_),
    .A2(_02525_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06888_ (.I(_01443_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06889_ (.A1(_02527_),
    .A2(_01451_),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06890_ (.A1(_01452_),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .B(_02528_),
    .C(\u_cpu.cpu.state.init_done ),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06891_ (.A1(_02520_),
    .A2(_02526_),
    .B1(_02529_),
    .B2(\u_cpu.cpu.state.stage_two_req ),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06892_ (.A1(\u_cpu.cpu.bufreg.lsb[0] ),
    .A2(_02530_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06893_ (.A1(_02524_),
    .A2(_02521_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06894_ (.A1(_02517_),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06895_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_02471_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06896_ (.A1(_02505_),
    .A2(_02469_),
    .A3(_02470_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06897_ (.A1(_02505_),
    .A2(_02534_),
    .B(_02535_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06898_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(\u_cpu.cpu.mem_bytecnt[0] ),
    .B(\u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06899_ (.A1(_02536_),
    .A2(_02537_),
    .B(_02533_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06900_ (.I(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06901_ (.A1(_01444_),
    .A2(_02463_),
    .B1(_02539_),
    .B2(_01460_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06902_ (.I(_02521_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06903_ (.I(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06904_ (.A1(_02541_),
    .A2(_02542_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06905_ (.A1(_02468_),
    .A2(_02540_),
    .A3(_02543_),
    .B(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06906_ (.I(_02544_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06907_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_02545_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06908_ (.A1(_02531_),
    .A2(_02533_),
    .B(_02538_),
    .C(_02546_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06909_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_02501_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06910_ (.A1(\u_cpu.cpu.bufreg.lsb[0] ),
    .A2(_02530_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06911_ (.A1(_02536_),
    .A2(_02537_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06912_ (.A1(_02533_),
    .A2(_02550_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06913_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_02544_),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06914_ (.A1(_02549_),
    .A2(_02533_),
    .B(_02551_),
    .C(_02552_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06915_ (.A1(_02547_),
    .A2(_02548_),
    .A3(_02553_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06916_ (.A1(_02518_),
    .A2(_02531_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06917_ (.A1(_02518_),
    .A2(_02554_),
    .B(_02555_),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06918_ (.I(_02527_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06919_ (.I(_02521_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06920_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_02478_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06921_ (.A1(_02485_),
    .A2(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06922_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_02478_),
    .B(_01452_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06923_ (.A1(_02492_),
    .A2(_02559_),
    .B(_02560_),
    .C(_02561_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06924_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .A3(_02479_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06925_ (.A1(_02485_),
    .A2(_02522_),
    .A3(\u_cpu.cpu.alu.cmp_r ),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06926_ (.A1(_01442_),
    .A2(_02563_),
    .B1(_02564_),
    .B2(_02548_),
    .C(_02549_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06927_ (.A1(_02562_),
    .A2(_02565_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06928_ (.A1(_02557_),
    .A2(_02518_),
    .A3(_02558_),
    .A4(_02566_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06929_ (.I(\u_cpu.cpu.mem_if.signbit ),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06930_ (.A1(_02491_),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .B1(\u_cpu.cpu.mem_bytecnt[0] ),
    .B2(_02486_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06931_ (.I0(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I3(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(\u_cpu.cpu.bufreg.lsb[0] ),
    .S1(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06932_ (.A1(_02569_),
    .A2(_02570_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06933_ (.A1(_02568_),
    .A2(_02569_),
    .B(_02571_),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06934_ (.A1(_02487_),
    .A2(_02571_),
    .B(_02524_),
    .C(_02558_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06935_ (.I(\u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06936_ (.A1(_02573_),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06937_ (.A1(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .B(_02500_),
    .C(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06938_ (.A1(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .A2(_02513_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06939_ (.A1(_02575_),
    .A2(_02576_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06940_ (.A1(_02517_),
    .A2(_02521_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06941_ (.A1(_02577_),
    .A2(_02578_),
    .B(_01463_),
    .C(_02510_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06942_ (.A1(_00798_),
    .A2(_02572_),
    .B(_02579_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06943_ (.A1(_02518_),
    .A2(_02532_),
    .A3(_02554_),
    .B(_02580_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06944_ (.A1(_02484_),
    .A2(_02556_),
    .B1(_02567_),
    .B2(_02581_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06945_ (.I(_02582_),
    .ZN(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06946_ (.I(\u_cpu.rf_ram_if.rtrig1 ),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06947_ (.I(_02583_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06948_ (.I(_02474_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06949_ (.A1(_02585_),
    .A2(\u_cpu.rf_ram.rdata[1] ),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06950_ (.I(_02583_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06951_ (.A1(_02587_),
    .A2(\u_cpu.rf_ram_if.rdata1[1] ),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06952_ (.A1(_02584_),
    .A2(_02586_),
    .B(_02588_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06953_ (.A1(_02585_),
    .A2(\u_cpu.rf_ram.rdata[2] ),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06954_ (.A1(_02587_),
    .A2(\u_cpu.rf_ram_if.rdata1[2] ),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06955_ (.A1(_02584_),
    .A2(_02589_),
    .B(_02590_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06956_ (.A1(_02585_),
    .A2(\u_cpu.rf_ram.rdata[3] ),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06957_ (.A1(_02587_),
    .A2(\u_cpu.rf_ram_if.rdata1[3] ),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06958_ (.A1(_02584_),
    .A2(_02591_),
    .B(_02592_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06959_ (.A1(_02474_),
    .A2(\u_cpu.rf_ram.rdata[4] ),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06960_ (.A1(_02583_),
    .A2(\u_cpu.rf_ram_if.rdata1[4] ),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06961_ (.A1(_02584_),
    .A2(_02593_),
    .B(_02594_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06962_ (.A1(_02474_),
    .A2(\u_cpu.rf_ram.rdata[5] ),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06963_ (.A1(_02583_),
    .A2(\u_cpu.rf_ram_if.rdata1[5] ),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06964_ (.A1(_02584_),
    .A2(_02595_),
    .B(_02596_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06965_ (.A1(_02474_),
    .A2(\u_cpu.rf_ram.rdata[6] ),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06966_ (.A1(_02583_),
    .A2(\u_cpu.rf_ram_if.rdata1[6] ),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06967_ (.A1(_02587_),
    .A2(_02597_),
    .B(_02598_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06968_ (.I(_01471_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06969_ (.A1(\u_cpu.rf_ram_if.rdata0[1] ),
    .A2(_02599_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06970_ (.A1(_01496_),
    .A2(_02475_),
    .B(_02600_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06971_ (.A1(\u_cpu.rf_ram_if.rdata0[2] ),
    .A2(_02599_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06972_ (.A1(_01496_),
    .A2(_02586_),
    .B(_02601_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06973_ (.I(_01471_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06974_ (.A1(\u_cpu.rf_ram_if.rdata0[3] ),
    .A2(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06975_ (.A1(_01496_),
    .A2(_02589_),
    .B(_02603_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06976_ (.A1(\u_cpu.rf_ram_if.rdata0[4] ),
    .A2(_02602_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06977_ (.A1(_01496_),
    .A2(_02591_),
    .B(_02604_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06978_ (.A1(\u_cpu.rf_ram_if.rdata0[5] ),
    .A2(_02602_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06979_ (.A1(_02599_),
    .A2(_02593_),
    .B(_02605_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06980_ (.A1(\u_cpu.rf_ram_if.rdata0[6] ),
    .A2(_02602_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06981_ (.A1(_02599_),
    .A2(_02595_),
    .B(_02606_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06982_ (.A1(\u_cpu.rf_ram_if.rdata0[7] ),
    .A2(_02602_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06983_ (.A1(_02599_),
    .A2(_02597_),
    .B(_02607_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06984_ (.I(net4),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06985_ (.I(_02608_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06986_ (.A1(net3),
    .A2(_02609_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06987_ (.I(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06988_ (.I(\u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06989_ (.A1(_02495_),
    .A2(_02611_),
    .B1(_02464_),
    .B2(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06990_ (.I(_02524_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06991_ (.I(_02518_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06992_ (.I(_02615_),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06993_ (.I(_02616_),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06994_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(_02498_),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06995_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_02618_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06996_ (.A1(_02614_),
    .A2(_02617_),
    .A3(_02619_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06997_ (.I(net2),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06998_ (.A1(_02621_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06999_ (.I(_02622_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07000_ (.A1(net4),
    .A2(_02623_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07001_ (.I(_02624_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07002_ (.A1(_02613_),
    .A2(_02620_),
    .B(_02625_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07003_ (.A1(_02610_),
    .A2(_02626_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07004_ (.I(_02463_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07005_ (.I(net4),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07006_ (.I(_02628_),
    .Z(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07007_ (.I(_02629_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07008_ (.A1(_02630_),
    .A2(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07009_ (.A1(_02627_),
    .A2(_02625_),
    .B(_02631_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07010_ (.I(\u_arbiter.i_wb_cpu_ack ),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07011_ (.I(_02608_),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07012_ (.I(_02633_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07013_ (.I(_02611_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07014_ (.A1(_02612_),
    .A2(_02635_),
    .B(_02633_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07015_ (.A1(_02632_),
    .A2(_02634_),
    .B(_02636_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07016_ (.I(_02637_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07017_ (.A1(_02492_),
    .A2(_02612_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07018_ (.A1(_02495_),
    .A2(_02629_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07019_ (.A1(_02611_),
    .A2(_02638_),
    .B(_02639_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07020_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_02634_),
    .B(_02640_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07021_ (.I(_02641_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07022_ (.I(\u_arbiter.i_wb_cpu_rdt[1] ),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07023_ (.I(_02629_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07024_ (.I(_02612_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07025_ (.A1(_02644_),
    .A2(_02635_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07026_ (.A1(_02642_),
    .A2(_02643_),
    .B1(_02645_),
    .B2(_02639_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07027_ (.I(\u_arbiter.i_wb_cpu_rdt[2] ),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07028_ (.A1(_02492_),
    .A2(_02612_),
    .B(_02635_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07029_ (.A1(_02646_),
    .A2(_02643_),
    .B1(_02639_),
    .B2(_02647_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07030_ (.I(\u_arbiter.i_wb_cpu_rdt[3] ),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07031_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07032_ (.A1(_02649_),
    .A2(_02609_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07033_ (.A1(_02648_),
    .A2(_02634_),
    .B(_02650_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07034_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07035_ (.I(_02633_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07036_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(_02651_),
    .S(_02652_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07037_ (.I(_02653_),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07038_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .S(_02652_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07039_ (.I(_02654_),
    .Z(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07040_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .S(_02652_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07041_ (.I(_02655_),
    .Z(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07042_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .S(_02652_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07043_ (.I(_02656_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07044_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .S(_02652_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07045_ (.I(_02657_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07046_ (.I(_02633_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07047_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .S(_02658_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07048_ (.I(_02659_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07049_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .S(_02658_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07050_ (.I(_02660_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07051_ (.I0(\u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .S(_02658_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07052_ (.I(_02661_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07053_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .S(_02658_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07054_ (.I(_02662_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07055_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .S(_02658_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07056_ (.I(_02663_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07057_ (.I(_02608_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07058_ (.I(_02664_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07059_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .S(_02665_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07060_ (.I(_02666_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07061_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .S(_02665_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07062_ (.I(_02667_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07063_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .S(_02665_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07064_ (.I(_02668_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07065_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .S(_02665_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07066_ (.I(_02669_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07067_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .S(_02665_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07068_ (.I(_02670_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07069_ (.I(_02664_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07070_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .S(_02671_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07071_ (.I(_02672_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07072_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .S(_02671_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07073_ (.I(_02673_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07074_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .S(_02671_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07075_ (.I(_02674_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07076_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .S(_02671_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07077_ (.I(_02675_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07078_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .S(_02671_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07079_ (.I(_02676_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07080_ (.I(_02664_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07081_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .S(_02677_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07082_ (.I(_02678_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07083_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .S(_02677_),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07084_ (.I(_02679_),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07085_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .S(_02677_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07086_ (.I(_02680_),
    .Z(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07087_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S(_02677_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07088_ (.I(_02681_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07089_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .S(_02677_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07090_ (.I(_02682_),
    .Z(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07091_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07092_ (.I(_02629_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07093_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_02684_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07094_ (.A1(_02683_),
    .A2(_02643_),
    .B(_02685_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07095_ (.I(_02664_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07096_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .S(_02686_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07097_ (.I(_02687_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07098_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .S(_02686_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07099_ (.I(_02688_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07100_ (.I0(\u_scanchain_local.module_data_in[34] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .S(_02686_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07101_ (.I(_02689_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07102_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07103_ (.A1(_02630_),
    .A2(\u_scanchain_local.module_data_in[35] ),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07104_ (.A1(_02690_),
    .A2(_02643_),
    .B(_02691_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07105_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07106_ (.A1(_02684_),
    .A2(\u_scanchain_local.module_data_in[36] ),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07107_ (.A1(_02692_),
    .A2(_02643_),
    .B(_02693_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07108_ (.A1(_02630_),
    .A2(\u_scanchain_local.module_data_in[37] ),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07109_ (.A1(_02628_),
    .A2(_02623_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07110_ (.I(_02695_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07111_ (.A1(_02513_),
    .A2(_02696_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07112_ (.A1(_02694_),
    .A2(_02697_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07113_ (.A1(_02630_),
    .A2(\u_scanchain_local.module_data_in[38] ),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07114_ (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07115_ (.A1(_02699_),
    .A2(_02696_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07116_ (.A1(_02698_),
    .A2(_02700_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07117_ (.I(_02608_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07118_ (.A1(_02621_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07119_ (.I(_02702_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07120_ (.A1(_02664_),
    .A2(_02703_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07121_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07122_ (.I(_02705_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07123_ (.I(_02706_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07124_ (.I(_02707_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07125_ (.I(_02708_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07126_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07127_ (.A1(_02709_),
    .A2(_02710_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _07128_ (.A1(_02701_),
    .A2(\u_scanchain_local.module_data_in[39] ),
    .B1(_02704_),
    .B2(_02711_),
    .C1(_02625_),
    .C2(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07129_ (.I(_02712_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07130_ (.I(_02695_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07131_ (.I(_02713_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07132_ (.I(_02709_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07133_ (.A1(_02715_),
    .A2(_02710_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07134_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_02716_),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07135_ (.A1(_02701_),
    .A2(\u_scanchain_local.module_data_in[40] ),
    .B1(_02625_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07136_ (.A1(_02714_),
    .A2(_02717_),
    .B(_02718_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07137_ (.A1(_02715_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(_02710_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07138_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_02719_),
    .Z(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07139_ (.I(_02608_),
    .Z(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07140_ (.I(_02624_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07141_ (.A1(_02721_),
    .A2(\u_scanchain_local.module_data_in[41] ),
    .B1(_02722_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07142_ (.A1(_02714_),
    .A2(_02720_),
    .B(_02723_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07143_ (.I(_02704_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07144_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07145_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _07146_ (.A1(_02726_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07147_ (.A1(_02725_),
    .A2(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07148_ (.A1(_02628_),
    .A2(_02702_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07149_ (.I(_02729_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07150_ (.A1(_02684_),
    .A2(\u_scanchain_local.module_data_in[42] ),
    .B1(_02730_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07151_ (.A1(_02724_),
    .A2(_02728_),
    .B(_02731_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07152_ (.A1(_02725_),
    .A2(_02727_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07153_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_02732_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07154_ (.A1(_02721_),
    .A2(\u_scanchain_local.module_data_in[43] ),
    .B1(_02722_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07155_ (.A1(_02714_),
    .A2(_02733_),
    .B(_02734_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07156_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_02725_),
    .A3(_02727_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07157_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_02735_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07158_ (.A1(_02721_),
    .A2(\u_scanchain_local.module_data_in[44] ),
    .B1(_02722_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07159_ (.A1(_02714_),
    .A2(_02736_),
    .B(_02737_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07160_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07161_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A4(_02727_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07162_ (.A1(_02738_),
    .A2(_02739_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07163_ (.A1(_02738_),
    .A2(_02739_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07164_ (.A1(_02696_),
    .A2(_02741_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07165_ (.A1(_02684_),
    .A2(\u_scanchain_local.module_data_in[45] ),
    .B1(_02730_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07166_ (.A1(_02740_),
    .A2(_02742_),
    .B(_02743_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07167_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07168_ (.A1(_02744_),
    .A2(_02738_),
    .A3(_02739_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07169_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_02740_),
    .B(_02713_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07170_ (.A1(_02684_),
    .A2(\u_scanchain_local.module_data_in[46] ),
    .B1(_02730_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07171_ (.A1(_02745_),
    .A2(_02746_),
    .B(_02747_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07172_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_02745_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07173_ (.I(_02628_),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07174_ (.A1(_02749_),
    .A2(\u_scanchain_local.module_data_in[47] ),
    .B1(_02730_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07175_ (.A1(_02724_),
    .A2(_02748_),
    .B(_02750_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07176_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07177_ (.A1(_02744_),
    .A2(_02738_),
    .A3(_02739_),
    .A4(_02751_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07178_ (.I(_02752_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07179_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_02745_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07180_ (.A1(_02753_),
    .A2(_02754_),
    .B(_02713_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07181_ (.A1(_02609_),
    .A2(\u_scanchain_local.module_data_in[48] ),
    .B1(_02625_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .C(_02755_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07182_ (.I(_02756_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07183_ (.I(_02623_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07184_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07185_ (.A1(_02758_),
    .A2(_02753_),
    .B(_02703_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07186_ (.A1(_02758_),
    .A2(_02753_),
    .B(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07187_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .A2(_02757_),
    .B(_02760_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07188_ (.A1(_02701_),
    .A2(\u_scanchain_local.module_data_in[49] ),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07189_ (.A1(_02634_),
    .A2(_02761_),
    .B(_02762_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07190_ (.I(_02704_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07191_ (.A1(_02758_),
    .A2(_02753_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07192_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_02753_),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07193_ (.I(_02629_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07194_ (.I(_02729_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07195_ (.A1(_02766_),
    .A2(\u_scanchain_local.module_data_in[50] ),
    .B1(_02767_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07196_ (.A1(_02763_),
    .A2(_02764_),
    .A3(_02765_),
    .B(_02768_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07197_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07198_ (.A1(_02769_),
    .A2(_02765_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07199_ (.A1(_02749_),
    .A2(\u_scanchain_local.module_data_in[51] ),
    .B1(_02730_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07200_ (.A1(_02724_),
    .A2(_02770_),
    .B(_02771_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07201_ (.A1(_02769_),
    .A2(_02765_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07202_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_02772_),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07203_ (.A1(_02721_),
    .A2(\u_scanchain_local.module_data_in[52] ),
    .B1(_02722_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07204_ (.A1(_02714_),
    .A2(_02773_),
    .B(_02774_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07205_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_02769_),
    .A3(_02765_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07206_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_02775_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07207_ (.A1(_02721_),
    .A2(\u_scanchain_local.module_data_in[53] ),
    .B1(_02722_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07208_ (.A1(_02696_),
    .A2(_02776_),
    .B(_02777_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07209_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07210_ (.A1(_02778_),
    .A2(_02775_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07211_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07212_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_02752_),
    .A4(_02780_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07213_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_02779_),
    .B(_02781_),
    .C(_02703_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07214_ (.I(_02623_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07215_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .A2(_02783_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07216_ (.A1(_02686_),
    .A2(_02782_),
    .A3(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07217_ (.A1(_02634_),
    .A2(\u_scanchain_local.module_data_in[54] ),
    .B(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07218_ (.I(_02786_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07219_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_02781_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07220_ (.I(_02729_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07221_ (.A1(_02749_),
    .A2(\u_scanchain_local.module_data_in[55] ),
    .B1(_02788_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07222_ (.A1(_02724_),
    .A2(_02787_),
    .B(_02789_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07223_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07224_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07225_ (.A1(_02790_),
    .A2(_02781_),
    .B(_02791_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07226_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A3(_02765_),
    .A4(_02780_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07227_ (.A1(_02703_),
    .A2(_02792_),
    .A3(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07228_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .A2(_02783_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07229_ (.A1(_02686_),
    .A2(_02794_),
    .A3(_02795_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07230_ (.A1(_02609_),
    .A2(\u_scanchain_local.module_data_in[56] ),
    .B(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07231_ (.I(_02797_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07232_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_02793_),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07233_ (.A1(_02749_),
    .A2(\u_scanchain_local.module_data_in[57] ),
    .B1(_02788_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07234_ (.A1(_02724_),
    .A2(_02798_),
    .B(_02799_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07235_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07236_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07237_ (.A1(_02801_),
    .A2(_02791_),
    .A3(_02790_),
    .A4(_02781_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07238_ (.A1(_02800_),
    .A2(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07239_ (.A1(_02800_),
    .A2(_02802_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07240_ (.A1(_02696_),
    .A2(_02804_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07241_ (.A1(_02749_),
    .A2(\u_scanchain_local.module_data_in[58] ),
    .B1(_02788_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07242_ (.A1(_02803_),
    .A2(_02805_),
    .B(_02806_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07243_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_02804_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07244_ (.I(_02628_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07245_ (.A1(_02808_),
    .A2(\u_scanchain_local.module_data_in[59] ),
    .B1(_02788_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07246_ (.A1(_02763_),
    .A2(_02807_),
    .B(_02809_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07247_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_02800_),
    .A3(_02802_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07248_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07249_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A4(_02802_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07250_ (.A1(_02703_),
    .A2(_02812_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07251_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .A2(_02783_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07252_ (.A1(_02811_),
    .A2(_02813_),
    .B(_02814_),
    .C(_02633_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07253_ (.A1(_02609_),
    .A2(\u_scanchain_local.module_data_in[60] ),
    .B(_02815_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07254_ (.I(_02816_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07255_ (.A1(_02701_),
    .A2(\u_scanchain_local.module_data_in[61] ),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07256_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A3(_02810_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07257_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07258_ (.A1(_02819_),
    .A2(_02812_),
    .B(_02783_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07259_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_02757_),
    .B1(_02818_),
    .B2(_02820_),
    .C(_02766_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07260_ (.A1(_02817_),
    .A2(_02821_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07261_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_02818_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07262_ (.A1(_02808_),
    .A2(\u_scanchain_local.module_data_in[62] ),
    .B1(_02788_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07263_ (.A1(_02763_),
    .A2(_02822_),
    .B(_02823_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07264_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07265_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07266_ (.A1(_02824_),
    .A2(_02825_),
    .A3(_02819_),
    .A4(_02812_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07267_ (.I(_02826_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07268_ (.A1(_02825_),
    .A2(_02818_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07269_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_02828_),
    .B(_02713_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07270_ (.A1(_02808_),
    .A2(\u_scanchain_local.module_data_in[63] ),
    .B1(_02767_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07271_ (.A1(_02827_),
    .A2(_02829_),
    .B(_02830_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07272_ (.I(\u_scanchain_local.module_data_in[64] ),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07273_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .Z(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07274_ (.A1(_02832_),
    .A2(_02827_),
    .B(_02783_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07275_ (.A1(_02832_),
    .A2(_02827_),
    .B(_02833_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07276_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_02757_),
    .B(_02766_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07277_ (.A1(_02630_),
    .A2(_02831_),
    .B1(_02834_),
    .B2(_02835_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07278_ (.A1(_02832_),
    .A2(_02827_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07279_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A3(_02827_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07280_ (.A1(_02713_),
    .A2(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07281_ (.A1(_02808_),
    .A2(\u_scanchain_local.module_data_in[65] ),
    .B1(_02767_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07282_ (.A1(_02836_),
    .A2(_02838_),
    .B(_02839_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07283_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_02837_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07284_ (.A1(_02808_),
    .A2(\u_scanchain_local.module_data_in[66] ),
    .B1(_02767_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07285_ (.A1(_02763_),
    .A2(_02840_),
    .B(_02841_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07286_ (.A1(_02701_),
    .A2(\u_scanchain_local.module_data_in[67] ),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07287_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A4(_02826_),
    .Z(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07288_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_02843_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07289_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_02843_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07290_ (.A1(_02757_),
    .A2(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07291_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_02757_),
    .B1(_02844_),
    .B2(_02846_),
    .C(_02766_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07292_ (.A1(_02842_),
    .A2(_02847_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07293_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_02844_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07294_ (.A1(_02766_),
    .A2(\u_scanchain_local.module_data_in[68] ),
    .B1(_02767_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07295_ (.A1(_02763_),
    .A2(_02848_),
    .B(_02849_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07296_ (.A1(_02615_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07297_ (.A1(_02615_),
    .A2(_02541_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07298_ (.A1(_02480_),
    .A2(\u_cpu.cpu.bufreg.c_r ),
    .A3(_02850_),
    .A4(_02851_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07299_ (.A1(_02558_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07300_ (.A1(_02853_),
    .A2(_02543_),
    .B(_02615_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07301_ (.A1(_02548_),
    .A2(_02854_),
    .B(_02557_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07302_ (.A1(_02536_),
    .A2(_02855_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07303_ (.A1(_02480_),
    .A2(_02850_),
    .A3(_02851_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07304_ (.A1(\u_cpu.cpu.bufreg.c_r ),
    .A2(_02857_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07305_ (.A1(_02856_),
    .A2(_02858_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07306_ (.A1(_02520_),
    .A2(_02526_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07307_ (.A1(\u_cpu.cpu.state.stage_two_req ),
    .A2(_02529_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07308_ (.A1(_02860_),
    .A2(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07309_ (.A1(_02852_),
    .A2(_02859_),
    .B(_02862_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07310_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_02545_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07311_ (.A1(_02519_),
    .A2(_02525_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07312_ (.A1(_02461_),
    .A2(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07313_ (.A1(_02863_),
    .A2(_02547_),
    .B(_02865_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07314_ (.A1(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .A2(_02513_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07315_ (.I(_02575_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07316_ (.A1(_02867_),
    .A2(_02576_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07317_ (.A1(_02866_),
    .A2(_02868_),
    .B(_02865_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07318_ (.I(_02618_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07319_ (.A1(_02484_),
    .A2(_01459_),
    .B(_02869_),
    .ZN(\u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07320_ (.I(\u_cpu.cpu.immdec.imm11_7[4] ),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07321_ (.I(\u_cpu.cpu.immdec.imm11_7[3] ),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _07322_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A3(_02871_),
    .A4(\u_cpu.cpu.immdec.imm11_7[0] ),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07323_ (.A1(_02558_),
    .A2(_02463_),
    .B(_02578_),
    .C(_02557_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07324_ (.I(_02864_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07325_ (.A1(_02870_),
    .A2(_02872_),
    .B(_02873_),
    .C(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07326_ (.A1(_02484_),
    .A2(_02875_),
    .B(_02869_),
    .ZN(\u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07327_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07328_ (.A1(_02514_),
    .A2(_01458_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07329_ (.A1(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .A2(_02514_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07330_ (.A1(_02876_),
    .A2(_02877_),
    .B1(_02878_),
    .B2(_02467_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07331_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_01449_),
    .A3(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07332_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07333_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_02881_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07334_ (.A1(_02484_),
    .A2(_02880_),
    .A3(_02882_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07335_ (.A1(_02879_),
    .A2(_02883_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07336_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07337_ (.A1(_02885_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .B(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07338_ (.A1(\u_cpu.raddr[0] ),
    .A2(_02886_),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07339_ (.I(_02887_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07340_ (.A1(_01591_),
    .A2(_02888_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07341_ (.A1(_02884_),
    .A2(_02889_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07342_ (.I(_02890_),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07343_ (.I(_02878_),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07344_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_02892_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07345_ (.I(\u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07346_ (.A1(_02876_),
    .A2(\u_cpu.rf_ram_if.wen1_r ),
    .B1(_01438_),
    .B2(\u_cpu.rf_ram_if.wen0_r ),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07347_ (.A1(_02894_),
    .A2(_02895_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07348_ (.A1(_02892_),
    .A2(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07349_ (.A1(_02871_),
    .A2(_02893_),
    .A3(_02897_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07350_ (.I(_02898_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07351_ (.A1(_02891_),
    .A2(_02899_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07352_ (.I(_02900_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07353_ (.I(_02881_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07354_ (.I(_02876_),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07355_ (.A1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .A2(_02903_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07356_ (.A1(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .A2(_02902_),
    .B(_02904_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07357_ (.I(_02905_),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07358_ (.I(_02906_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07359_ (.I(_02907_),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07360_ (.I(_02900_),
    .Z(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07361_ (.A1(\u_cpu.rf_ram.memory[82][0] ),
    .A2(_02909_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07362_ (.A1(_02901_),
    .A2(_02908_),
    .B(_02910_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07363_ (.A1(_02903_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .Z(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07364_ (.A1(_02902_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .B(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07365_ (.I(_02912_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07366_ (.I(_02913_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07367_ (.I(_02914_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07368_ (.A1(\u_cpu.rf_ram.memory[82][1] ),
    .A2(_02909_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07369_ (.A1(_02901_),
    .A2(_02915_),
    .B(_02916_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07370_ (.A1(_02903_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .Z(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07371_ (.A1(_02902_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .B(_02917_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07372_ (.I(_02918_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07373_ (.I(_02919_),
    .Z(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07374_ (.I(_02920_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07375_ (.I(_02900_),
    .Z(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07376_ (.A1(\u_cpu.rf_ram.memory[82][2] ),
    .A2(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07377_ (.A1(_02901_),
    .A2(_02921_),
    .B(_02923_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07378_ (.A1(_02903_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07379_ (.A1(_02902_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .B(_02924_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07380_ (.I(_02925_),
    .Z(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07381_ (.I(_02926_),
    .Z(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07382_ (.I(_02927_),
    .Z(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07383_ (.A1(\u_cpu.rf_ram.memory[82][3] ),
    .A2(_02922_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07384_ (.A1(_02901_),
    .A2(_02928_),
    .B(_02929_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07385_ (.A1(_02903_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .Z(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07386_ (.A1(_02902_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .B(_02930_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07387_ (.I(_02931_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07388_ (.I(_02932_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07389_ (.I(_02933_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07390_ (.A1(\u_cpu.rf_ram.memory[82][4] ),
    .A2(_02922_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07391_ (.A1(_02901_),
    .A2(_02934_),
    .B(_02935_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07392_ (.A1(_02876_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07393_ (.A1(_02881_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .B(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07394_ (.I(_02937_),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07395_ (.I(_02938_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07396_ (.I(_02939_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07397_ (.A1(\u_cpu.rf_ram.memory[82][5] ),
    .A2(_02922_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07398_ (.A1(_02909_),
    .A2(_02940_),
    .B(_02941_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07399_ (.A1(_02876_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07400_ (.A1(_02881_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .B(_02942_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07401_ (.I(_02943_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07402_ (.I(_02944_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07403_ (.I(_02945_),
    .Z(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07404_ (.A1(\u_cpu.rf_ram.memory[82][6] ),
    .A2(_02922_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07405_ (.A1(_02909_),
    .A2(_02946_),
    .B(_02947_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07406_ (.I(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07407_ (.I0(_02948_),
    .I1(_02582_),
    .S(_02881_),
    .Z(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07408_ (.I(_02949_),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07409_ (.I(_02950_),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07410_ (.I(_02951_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07411_ (.A1(\u_cpu.rf_ram.memory[82][7] ),
    .A2(_02900_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07412_ (.A1(_02909_),
    .A2(_02952_),
    .B(_02953_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07413_ (.I(_02906_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07414_ (.A1(_02885_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .B(\u_cpu.raddr[0] ),
    .C(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07415_ (.A1(\u_cpu.raddr[1] ),
    .A2(_02955_),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07416_ (.A1(_02888_),
    .A2(_02956_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07417_ (.A1(_01463_),
    .A2(_02880_),
    .A3(_02882_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07418_ (.A1(_02879_),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07419_ (.A1(_02957_),
    .A2(_02959_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07420_ (.I(_02960_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07421_ (.I(_02895_),
    .Z(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07422_ (.A1(_02871_),
    .A2(_02870_),
    .A3(_02893_),
    .A4(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07423_ (.I(_02963_),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07424_ (.A1(_02961_),
    .A2(_02964_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07425_ (.I(_02965_),
    .Z(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07426_ (.I(_02965_),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07427_ (.A1(\u_cpu.rf_ram.memory[21][0] ),
    .A2(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07428_ (.A1(_02954_),
    .A2(_02966_),
    .B(_02968_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07429_ (.I(_02913_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07430_ (.A1(\u_cpu.rf_ram.memory[21][1] ),
    .A2(_02967_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07431_ (.A1(_02969_),
    .A2(_02966_),
    .B(_02970_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07432_ (.I(_02919_),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07433_ (.I(_02965_),
    .Z(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07434_ (.A1(\u_cpu.rf_ram.memory[21][2] ),
    .A2(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07435_ (.A1(_02971_),
    .A2(_02966_),
    .B(_02973_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07436_ (.I(_02926_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07437_ (.A1(\u_cpu.rf_ram.memory[21][3] ),
    .A2(_02972_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07438_ (.A1(_02974_),
    .A2(_02966_),
    .B(_02975_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07439_ (.I(_02932_),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07440_ (.A1(\u_cpu.rf_ram.memory[21][4] ),
    .A2(_02972_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07441_ (.A1(_02976_),
    .A2(_02966_),
    .B(_02977_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07442_ (.I(_02938_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07443_ (.A1(\u_cpu.rf_ram.memory[21][5] ),
    .A2(_02972_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07444_ (.A1(_02978_),
    .A2(_02967_),
    .B(_02979_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07445_ (.I(_02944_),
    .Z(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07446_ (.A1(\u_cpu.rf_ram.memory[21][6] ),
    .A2(_02972_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07447_ (.A1(_02980_),
    .A2(_02967_),
    .B(_02981_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07448_ (.I(_02950_),
    .Z(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07449_ (.A1(\u_cpu.rf_ram.memory[21][7] ),
    .A2(_02965_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07450_ (.A1(_02982_),
    .A2(_02967_),
    .B(_02983_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07451_ (.A1(_02884_),
    .A2(_02957_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07452_ (.I(_02984_),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07453_ (.A1(_02899_),
    .A2(_02985_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07454_ (.I(_02986_),
    .Z(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07455_ (.I(_02986_),
    .Z(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07456_ (.A1(\u_cpu.rf_ram.memory[81][0] ),
    .A2(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07457_ (.A1(_02954_),
    .A2(_02987_),
    .B(_02989_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07458_ (.A1(\u_cpu.rf_ram.memory[81][1] ),
    .A2(_02988_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07459_ (.A1(_02969_),
    .A2(_02987_),
    .B(_02990_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07460_ (.I(_02986_),
    .Z(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07461_ (.A1(\u_cpu.rf_ram.memory[81][2] ),
    .A2(_02991_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07462_ (.A1(_02971_),
    .A2(_02987_),
    .B(_02992_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07463_ (.A1(\u_cpu.rf_ram.memory[81][3] ),
    .A2(_02991_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07464_ (.A1(_02974_),
    .A2(_02987_),
    .B(_02993_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07465_ (.A1(\u_cpu.rf_ram.memory[81][4] ),
    .A2(_02991_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07466_ (.A1(_02976_),
    .A2(_02987_),
    .B(_02994_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07467_ (.A1(\u_cpu.rf_ram.memory[81][5] ),
    .A2(_02991_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07468_ (.A1(_02978_),
    .A2(_02988_),
    .B(_02995_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07469_ (.A1(\u_cpu.rf_ram.memory[81][6] ),
    .A2(_02991_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07470_ (.A1(_02980_),
    .A2(_02988_),
    .B(_02996_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07471_ (.A1(\u_cpu.rf_ram.memory[81][7] ),
    .A2(_02986_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07472_ (.A1(_02982_),
    .A2(_02988_),
    .B(_02997_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07473_ (.A1(_02891_),
    .A2(_02964_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07474_ (.I(_02998_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07475_ (.I(_02998_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07476_ (.A1(\u_cpu.rf_ram.memory[18][0] ),
    .A2(_03000_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07477_ (.A1(_02954_),
    .A2(_02999_),
    .B(_03001_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07478_ (.A1(\u_cpu.rf_ram.memory[18][1] ),
    .A2(_03000_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07479_ (.A1(_02969_),
    .A2(_02999_),
    .B(_03002_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07480_ (.I(_02998_),
    .Z(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07481_ (.A1(\u_cpu.rf_ram.memory[18][2] ),
    .A2(_03003_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07482_ (.A1(_02971_),
    .A2(_02999_),
    .B(_03004_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07483_ (.A1(\u_cpu.rf_ram.memory[18][3] ),
    .A2(_03003_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07484_ (.A1(_02974_),
    .A2(_02999_),
    .B(_03005_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07485_ (.A1(\u_cpu.rf_ram.memory[18][4] ),
    .A2(_03003_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07486_ (.A1(_02976_),
    .A2(_02999_),
    .B(_03006_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07487_ (.A1(\u_cpu.rf_ram.memory[18][5] ),
    .A2(_03003_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07488_ (.A1(_02978_),
    .A2(_03000_),
    .B(_03007_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07489_ (.A1(\u_cpu.rf_ram.memory[18][6] ),
    .A2(_03003_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07490_ (.A1(_02980_),
    .A2(_03000_),
    .B(_03008_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07491_ (.A1(\u_cpu.rf_ram.memory[18][7] ),
    .A2(_02998_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07492_ (.A1(_02982_),
    .A2(_03000_),
    .B(_03009_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07493_ (.I(_02907_),
    .Z(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07494_ (.A1(_01591_),
    .A2(_02887_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07495_ (.A1(_02959_),
    .A2(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07496_ (.I(_03012_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07497_ (.A1(_02964_),
    .A2(_03013_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07498_ (.I(_03014_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07499_ (.I(_03014_),
    .Z(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07500_ (.A1(\u_cpu.rf_ram.memory[20][0] ),
    .A2(_03016_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07501_ (.A1(_03010_),
    .A2(_03015_),
    .B(_03017_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07502_ (.I(_02914_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07503_ (.A1(\u_cpu.rf_ram.memory[20][1] ),
    .A2(_03016_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07504_ (.A1(_03018_),
    .A2(_03015_),
    .B(_03019_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07505_ (.I(_02920_),
    .Z(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07506_ (.I(_03014_),
    .Z(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07507_ (.A1(\u_cpu.rf_ram.memory[20][2] ),
    .A2(_03021_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07508_ (.A1(_03020_),
    .A2(_03015_),
    .B(_03022_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07509_ (.I(_02927_),
    .Z(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07510_ (.A1(\u_cpu.rf_ram.memory[20][3] ),
    .A2(_03021_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07511_ (.A1(_03023_),
    .A2(_03015_),
    .B(_03024_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07512_ (.I(_02933_),
    .Z(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07513_ (.A1(\u_cpu.rf_ram.memory[20][4] ),
    .A2(_03021_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07514_ (.A1(_03025_),
    .A2(_03015_),
    .B(_03026_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07515_ (.I(_02939_),
    .Z(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07516_ (.A1(\u_cpu.rf_ram.memory[20][5] ),
    .A2(_03021_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07517_ (.A1(_03027_),
    .A2(_03016_),
    .B(_03028_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07518_ (.I(_02945_),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07519_ (.A1(\u_cpu.rf_ram.memory[20][6] ),
    .A2(_03021_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07520_ (.A1(_03029_),
    .A2(_03016_),
    .B(_03030_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07521_ (.I(_02951_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07522_ (.A1(\u_cpu.rf_ram.memory[20][7] ),
    .A2(_03014_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07523_ (.A1(_03031_),
    .A2(_03016_),
    .B(_03032_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07524_ (.I(\u_cpu.cpu.immdec.imm11_7[2] ),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07525_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_02878_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07526_ (.A1(_03033_),
    .A2(_02892_),
    .A3(_03034_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07527_ (.A1(_02870_),
    .A2(_02962_),
    .A3(_03035_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07528_ (.I(_03036_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07529_ (.A1(_02985_),
    .A2(_03037_),
    .Z(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07530_ (.I(_03038_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07531_ (.I(_03038_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07532_ (.A1(\u_cpu.rf_ram.memory[1][0] ),
    .A2(_03040_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07533_ (.A1(_02908_),
    .A2(_03039_),
    .B(_03041_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07534_ (.A1(\u_cpu.rf_ram.memory[1][1] ),
    .A2(_03040_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07535_ (.A1(_02915_),
    .A2(_03039_),
    .B(_03042_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07536_ (.I(_03038_),
    .Z(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07537_ (.A1(\u_cpu.rf_ram.memory[1][2] ),
    .A2(_03043_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07538_ (.A1(_02921_),
    .A2(_03039_),
    .B(_03044_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07539_ (.A1(\u_cpu.rf_ram.memory[1][3] ),
    .A2(_03043_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07540_ (.A1(_02928_),
    .A2(_03039_),
    .B(_03045_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07541_ (.A1(\u_cpu.rf_ram.memory[1][4] ),
    .A2(_03043_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07542_ (.A1(_02934_),
    .A2(_03039_),
    .B(_03046_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07543_ (.A1(\u_cpu.rf_ram.memory[1][5] ),
    .A2(_03043_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07544_ (.A1(_02940_),
    .A2(_03040_),
    .B(_03047_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07545_ (.A1(\u_cpu.rf_ram.memory[1][6] ),
    .A2(_03043_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07546_ (.A1(_02946_),
    .A2(_03040_),
    .B(_03048_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07547_ (.A1(\u_cpu.rf_ram.memory[1][7] ),
    .A2(_03038_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07548_ (.A1(_02952_),
    .A2(_03040_),
    .B(_03049_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07549_ (.I(_03036_),
    .Z(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07550_ (.A1(_02887_),
    .A2(_02956_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07551_ (.A1(_02959_),
    .A2(_03051_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07552_ (.I(_03052_),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07553_ (.A1(_03050_),
    .A2(_03053_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07554_ (.I(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07555_ (.I(_03055_),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07556_ (.I(_03055_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07557_ (.A1(\u_cpu.rf_ram.memory[7][0] ),
    .A2(_03057_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07558_ (.A1(_02908_),
    .A2(_03056_),
    .B(_03058_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07559_ (.A1(\u_cpu.rf_ram.memory[7][1] ),
    .A2(_03057_),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07560_ (.A1(_02915_),
    .A2(_03056_),
    .B(_03059_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07561_ (.I(_03055_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07562_ (.A1(\u_cpu.rf_ram.memory[7][2] ),
    .A2(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07563_ (.A1(_02921_),
    .A2(_03056_),
    .B(_03061_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07564_ (.A1(\u_cpu.rf_ram.memory[7][3] ),
    .A2(_03060_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07565_ (.A1(_02928_),
    .A2(_03056_),
    .B(_03062_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07566_ (.A1(\u_cpu.rf_ram.memory[7][4] ),
    .A2(_03060_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07567_ (.A1(_02934_),
    .A2(_03056_),
    .B(_03063_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07568_ (.A1(\u_cpu.rf_ram.memory[7][5] ),
    .A2(_03060_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07569_ (.A1(_02940_),
    .A2(_03057_),
    .B(_03064_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07570_ (.A1(\u_cpu.rf_ram.memory[7][6] ),
    .A2(_03060_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07571_ (.A1(_02946_),
    .A2(_03057_),
    .B(_03065_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07572_ (.A1(\u_cpu.rf_ram.memory[7][7] ),
    .A2(_03055_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07573_ (.A1(_02952_),
    .A2(_03057_),
    .B(_03066_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07574_ (.A1(_02884_),
    .A2(_03011_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07575_ (.I(_03067_),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07576_ (.A1(_02899_),
    .A2(_03068_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07577_ (.I(_03069_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07578_ (.I(_03069_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07579_ (.A1(\u_cpu.rf_ram.memory[80][0] ),
    .A2(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07580_ (.A1(_03010_),
    .A2(_03070_),
    .B(_03072_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07581_ (.A1(\u_cpu.rf_ram.memory[80][1] ),
    .A2(_03071_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07582_ (.A1(_03018_),
    .A2(_03070_),
    .B(_03073_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07583_ (.I(_03069_),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07584_ (.A1(\u_cpu.rf_ram.memory[80][2] ),
    .A2(_03074_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07585_ (.A1(_03020_),
    .A2(_03070_),
    .B(_03075_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07586_ (.A1(\u_cpu.rf_ram.memory[80][3] ),
    .A2(_03074_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07587_ (.A1(_03023_),
    .A2(_03070_),
    .B(_03076_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07588_ (.A1(\u_cpu.rf_ram.memory[80][4] ),
    .A2(_03074_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07589_ (.A1(_03025_),
    .A2(_03070_),
    .B(_03077_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07590_ (.A1(\u_cpu.rf_ram.memory[80][5] ),
    .A2(_03074_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07591_ (.A1(_03027_),
    .A2(_03071_),
    .B(_03078_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07592_ (.A1(\u_cpu.rf_ram.memory[80][6] ),
    .A2(_03074_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07593_ (.A1(_03029_),
    .A2(_03071_),
    .B(_03079_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07594_ (.A1(\u_cpu.rf_ram.memory[80][7] ),
    .A2(_03069_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07595_ (.A1(_03031_),
    .A2(_03071_),
    .B(_03080_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07596_ (.A1(_02879_),
    .A2(_02883_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07597_ (.A1(_02889_),
    .A2(_03081_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07598_ (.I(_03082_),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07599_ (.I(_03033_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07600_ (.I(_03034_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07601_ (.A1(_03084_),
    .A2(_02892_),
    .A3(_02896_),
    .A4(_03085_),
    .Z(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07602_ (.I(_03086_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07603_ (.A1(_03083_),
    .A2(_03087_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07604_ (.I(_03088_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07605_ (.I(_03088_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07606_ (.A1(\u_cpu.rf_ram.memory[78][0] ),
    .A2(_03090_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07607_ (.A1(_03010_),
    .A2(_03089_),
    .B(_03091_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07608_ (.A1(\u_cpu.rf_ram.memory[78][1] ),
    .A2(_03090_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07609_ (.A1(_03018_),
    .A2(_03089_),
    .B(_03092_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07610_ (.I(_03088_),
    .Z(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07611_ (.A1(\u_cpu.rf_ram.memory[78][2] ),
    .A2(_03093_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07612_ (.A1(_03020_),
    .A2(_03089_),
    .B(_03094_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07613_ (.A1(\u_cpu.rf_ram.memory[78][3] ),
    .A2(_03093_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07614_ (.A1(_03023_),
    .A2(_03089_),
    .B(_03095_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07615_ (.A1(\u_cpu.rf_ram.memory[78][4] ),
    .A2(_03093_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07616_ (.A1(_03025_),
    .A2(_03089_),
    .B(_03096_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07617_ (.A1(\u_cpu.rf_ram.memory[78][5] ),
    .A2(_03093_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07618_ (.A1(_03027_),
    .A2(_03090_),
    .B(_03097_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07619_ (.A1(\u_cpu.rf_ram.memory[78][6] ),
    .A2(_03093_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07620_ (.A1(_03029_),
    .A2(_03090_),
    .B(_03098_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07621_ (.A1(\u_cpu.rf_ram.memory[78][7] ),
    .A2(_03088_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07622_ (.A1(_03031_),
    .A2(_03090_),
    .B(_03099_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07623_ (.A1(_02879_),
    .A2(_02958_),
    .Z(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07624_ (.A1(_02889_),
    .A2(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07625_ (.I(_03101_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07626_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A3(_02962_),
    .A4(_03085_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07627_ (.I(_03103_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07628_ (.A1(_03102_),
    .A2(_03104_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07629_ (.I(_03105_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07630_ (.I(_03105_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07631_ (.A1(\u_cpu.rf_ram.memory[42][0] ),
    .A2(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07632_ (.A1(_03010_),
    .A2(_03106_),
    .B(_03108_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07633_ (.A1(\u_cpu.rf_ram.memory[42][1] ),
    .A2(_03107_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07634_ (.A1(_03018_),
    .A2(_03106_),
    .B(_03109_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07635_ (.I(_03105_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07636_ (.A1(\u_cpu.rf_ram.memory[42][2] ),
    .A2(_03110_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07637_ (.A1(_03020_),
    .A2(_03106_),
    .B(_03111_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07638_ (.A1(\u_cpu.rf_ram.memory[42][3] ),
    .A2(_03110_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07639_ (.A1(_03023_),
    .A2(_03106_),
    .B(_03112_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07640_ (.A1(\u_cpu.rf_ram.memory[42][4] ),
    .A2(_03110_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07641_ (.A1(_03025_),
    .A2(_03106_),
    .B(_03113_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07642_ (.A1(\u_cpu.rf_ram.memory[42][5] ),
    .A2(_03110_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07643_ (.A1(_03027_),
    .A2(_03107_),
    .B(_03114_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07644_ (.A1(\u_cpu.rf_ram.memory[42][6] ),
    .A2(_03110_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07645_ (.A1(_03029_),
    .A2(_03107_),
    .B(_03115_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07646_ (.A1(\u_cpu.rf_ram.memory[42][7] ),
    .A2(_03105_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07647_ (.A1(_03031_),
    .A2(_03107_),
    .B(_03116_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07648_ (.A1(_03083_),
    .A2(_03104_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07649_ (.I(_03117_),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07650_ (.I(_03117_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07651_ (.A1(\u_cpu.rf_ram.memory[46][0] ),
    .A2(_03119_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07652_ (.A1(_03010_),
    .A2(_03118_),
    .B(_03120_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07653_ (.A1(\u_cpu.rf_ram.memory[46][1] ),
    .A2(_03119_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07654_ (.A1(_03018_),
    .A2(_03118_),
    .B(_03121_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07655_ (.I(_03117_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07656_ (.A1(\u_cpu.rf_ram.memory[46][2] ),
    .A2(_03122_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07657_ (.A1(_03020_),
    .A2(_03118_),
    .B(_03123_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07658_ (.A1(\u_cpu.rf_ram.memory[46][3] ),
    .A2(_03122_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07659_ (.A1(_03023_),
    .A2(_03118_),
    .B(_03124_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07660_ (.A1(\u_cpu.rf_ram.memory[46][4] ),
    .A2(_03122_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07661_ (.A1(_03025_),
    .A2(_03118_),
    .B(_03125_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07662_ (.A1(\u_cpu.rf_ram.memory[46][5] ),
    .A2(_03122_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07663_ (.A1(_03027_),
    .A2(_03119_),
    .B(_03126_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07664_ (.A1(\u_cpu.rf_ram.memory[46][6] ),
    .A2(_03122_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07665_ (.A1(_03029_),
    .A2(_03119_),
    .B(_03127_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07666_ (.A1(\u_cpu.rf_ram.memory[46][7] ),
    .A2(_03117_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07667_ (.A1(_03031_),
    .A2(_03119_),
    .B(_03128_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07668_ (.I(_02907_),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07669_ (.I(_03103_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07670_ (.A1(_02957_),
    .A2(_03081_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07671_ (.I(_03131_),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07672_ (.A1(_03130_),
    .A2(_03132_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07673_ (.I(_03133_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07674_ (.I(_03133_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07675_ (.A1(\u_cpu.rf_ram.memory[45][0] ),
    .A2(_03135_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07676_ (.A1(_03129_),
    .A2(_03134_),
    .B(_03136_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07677_ (.I(_02914_),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07678_ (.A1(\u_cpu.rf_ram.memory[45][1] ),
    .A2(_03135_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07679_ (.A1(_03137_),
    .A2(_03134_),
    .B(_03138_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07680_ (.I(_02920_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07681_ (.I(_03133_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07682_ (.A1(\u_cpu.rf_ram.memory[45][2] ),
    .A2(_03140_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07683_ (.A1(_03139_),
    .A2(_03134_),
    .B(_03141_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07684_ (.I(_02927_),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07685_ (.A1(\u_cpu.rf_ram.memory[45][3] ),
    .A2(_03140_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07686_ (.A1(_03142_),
    .A2(_03134_),
    .B(_03143_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07687_ (.I(_02933_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07688_ (.A1(\u_cpu.rf_ram.memory[45][4] ),
    .A2(_03140_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07689_ (.A1(_03144_),
    .A2(_03134_),
    .B(_03145_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07690_ (.I(_02939_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07691_ (.A1(\u_cpu.rf_ram.memory[45][5] ),
    .A2(_03140_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07692_ (.A1(_03146_),
    .A2(_03135_),
    .B(_03147_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07693_ (.I(_02945_),
    .Z(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07694_ (.A1(\u_cpu.rf_ram.memory[45][6] ),
    .A2(_03140_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07695_ (.A1(_03148_),
    .A2(_03135_),
    .B(_03149_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07696_ (.I(_02951_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07697_ (.A1(\u_cpu.rf_ram.memory[45][7] ),
    .A2(_03133_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07698_ (.A1(_03150_),
    .A2(_03135_),
    .B(_03151_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07699_ (.A1(_03011_),
    .A2(_03081_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07700_ (.I(_03152_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07701_ (.A1(_03130_),
    .A2(_03153_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07702_ (.I(_03154_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07703_ (.I(_03154_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07704_ (.A1(\u_cpu.rf_ram.memory[44][0] ),
    .A2(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07705_ (.A1(_03129_),
    .A2(_03155_),
    .B(_03157_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07706_ (.A1(\u_cpu.rf_ram.memory[44][1] ),
    .A2(_03156_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07707_ (.A1(_03137_),
    .A2(_03155_),
    .B(_03158_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07708_ (.I(_03154_),
    .Z(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07709_ (.A1(\u_cpu.rf_ram.memory[44][2] ),
    .A2(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07710_ (.A1(_03139_),
    .A2(_03155_),
    .B(_03160_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07711_ (.A1(\u_cpu.rf_ram.memory[44][3] ),
    .A2(_03159_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07712_ (.A1(_03142_),
    .A2(_03155_),
    .B(_03161_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07713_ (.A1(\u_cpu.rf_ram.memory[44][4] ),
    .A2(_03159_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07714_ (.A1(_03144_),
    .A2(_03155_),
    .B(_03162_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07715_ (.A1(\u_cpu.rf_ram.memory[44][5] ),
    .A2(_03159_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07716_ (.A1(_03146_),
    .A2(_03156_),
    .B(_03163_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07717_ (.A1(\u_cpu.rf_ram.memory[44][6] ),
    .A2(_03159_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07718_ (.A1(_03148_),
    .A2(_03156_),
    .B(_03164_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07719_ (.A1(\u_cpu.rf_ram.memory[44][7] ),
    .A2(_03154_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07720_ (.A1(_03150_),
    .A2(_03156_),
    .B(_03165_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07721_ (.A1(_02884_),
    .A2(_03051_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07722_ (.A1(_03084_),
    .A2(_02870_),
    .A3(_02962_),
    .A4(_03085_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07723_ (.I(_03167_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07724_ (.A1(_03166_),
    .A2(_03168_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07725_ (.I(_03169_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07726_ (.I(_03169_),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07727_ (.A1(\u_cpu.rf_ram.memory[51][0] ),
    .A2(_03171_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07728_ (.A1(_03129_),
    .A2(_03170_),
    .B(_03172_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07729_ (.A1(\u_cpu.rf_ram.memory[51][1] ),
    .A2(_03171_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07730_ (.A1(_03137_),
    .A2(_03170_),
    .B(_03173_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07731_ (.I(_03169_),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07732_ (.A1(\u_cpu.rf_ram.memory[51][2] ),
    .A2(_03174_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07733_ (.A1(_03139_),
    .A2(_03170_),
    .B(_03175_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07734_ (.A1(\u_cpu.rf_ram.memory[51][3] ),
    .A2(_03174_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07735_ (.A1(_03142_),
    .A2(_03170_),
    .B(_03176_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07736_ (.A1(\u_cpu.rf_ram.memory[51][4] ),
    .A2(_03174_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07737_ (.A1(_03144_),
    .A2(_03170_),
    .B(_03177_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07738_ (.A1(\u_cpu.rf_ram.memory[51][5] ),
    .A2(_03174_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07739_ (.A1(_03146_),
    .A2(_03171_),
    .B(_03178_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07740_ (.A1(\u_cpu.rf_ram.memory[51][6] ),
    .A2(_03174_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07741_ (.A1(_03148_),
    .A2(_03171_),
    .B(_03179_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07742_ (.A1(\u_cpu.rf_ram.memory[51][7] ),
    .A2(_03169_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07743_ (.A1(_03150_),
    .A2(_03171_),
    .B(_03180_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07744_ (.I(_03103_),
    .Z(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07745_ (.A1(_02957_),
    .A2(_03100_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07746_ (.I(_03182_),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07747_ (.A1(_03181_),
    .A2(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07748_ (.I(_03184_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07749_ (.I(_03184_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07750_ (.A1(\u_cpu.rf_ram.memory[41][0] ),
    .A2(_03186_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07751_ (.A1(_03129_),
    .A2(_03185_),
    .B(_03187_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07752_ (.A1(\u_cpu.rf_ram.memory[41][1] ),
    .A2(_03186_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07753_ (.A1(_03137_),
    .A2(_03185_),
    .B(_03188_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07754_ (.I(_03184_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07755_ (.A1(\u_cpu.rf_ram.memory[41][2] ),
    .A2(_03189_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07756_ (.A1(_03139_),
    .A2(_03185_),
    .B(_03190_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07757_ (.A1(\u_cpu.rf_ram.memory[41][3] ),
    .A2(_03189_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07758_ (.A1(_03142_),
    .A2(_03185_),
    .B(_03191_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07759_ (.A1(\u_cpu.rf_ram.memory[41][4] ),
    .A2(_03189_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07760_ (.A1(_03144_),
    .A2(_03185_),
    .B(_03192_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07761_ (.A1(\u_cpu.rf_ram.memory[41][5] ),
    .A2(_03189_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07762_ (.A1(_03146_),
    .A2(_03186_),
    .B(_03193_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07763_ (.A1(\u_cpu.rf_ram.memory[41][6] ),
    .A2(_03189_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07764_ (.A1(_03148_),
    .A2(_03186_),
    .B(_03194_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07765_ (.A1(\u_cpu.rf_ram.memory[41][7] ),
    .A2(_03184_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07766_ (.A1(_03150_),
    .A2(_03186_),
    .B(_03195_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07767_ (.A1(_03051_),
    .A2(_03100_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07768_ (.I(_03196_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07769_ (.A1(_03181_),
    .A2(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07770_ (.I(_03198_),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07771_ (.I(_03198_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07772_ (.A1(\u_cpu.rf_ram.memory[43][0] ),
    .A2(_03200_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07773_ (.A1(_03129_),
    .A2(_03199_),
    .B(_03201_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07774_ (.A1(\u_cpu.rf_ram.memory[43][1] ),
    .A2(_03200_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07775_ (.A1(_03137_),
    .A2(_03199_),
    .B(_03202_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07776_ (.I(_03198_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07777_ (.A1(\u_cpu.rf_ram.memory[43][2] ),
    .A2(_03203_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07778_ (.A1(_03139_),
    .A2(_03199_),
    .B(_03204_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07779_ (.A1(\u_cpu.rf_ram.memory[43][3] ),
    .A2(_03203_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07780_ (.A1(_03142_),
    .A2(_03199_),
    .B(_03205_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07781_ (.A1(\u_cpu.rf_ram.memory[43][4] ),
    .A2(_03203_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07782_ (.A1(_03144_),
    .A2(_03199_),
    .B(_03206_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07783_ (.A1(\u_cpu.rf_ram.memory[43][5] ),
    .A2(_03203_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07784_ (.A1(_03146_),
    .A2(_03200_),
    .B(_03207_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07785_ (.A1(\u_cpu.rf_ram.memory[43][6] ),
    .A2(_03203_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07786_ (.A1(_03148_),
    .A2(_03200_),
    .B(_03208_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07787_ (.A1(\u_cpu.rf_ram.memory[43][7] ),
    .A2(_03198_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07788_ (.A1(_03150_),
    .A2(_03200_),
    .B(_03209_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07789_ (.I(_02907_),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07790_ (.A1(_03068_),
    .A2(_03168_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07791_ (.I(_03211_),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07792_ (.I(_03211_),
    .Z(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07793_ (.A1(\u_cpu.rf_ram.memory[48][0] ),
    .A2(_03213_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07794_ (.A1(_03210_),
    .A2(_03212_),
    .B(_03214_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07795_ (.I(_02914_),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07796_ (.A1(\u_cpu.rf_ram.memory[48][1] ),
    .A2(_03213_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07797_ (.A1(_03215_),
    .A2(_03212_),
    .B(_03216_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07798_ (.I(_02920_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07799_ (.I(_03211_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07800_ (.A1(\u_cpu.rf_ram.memory[48][2] ),
    .A2(_03218_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07801_ (.A1(_03217_),
    .A2(_03212_),
    .B(_03219_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07802_ (.I(_02927_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07803_ (.A1(\u_cpu.rf_ram.memory[48][3] ),
    .A2(_03218_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07804_ (.A1(_03220_),
    .A2(_03212_),
    .B(_03221_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07805_ (.I(_02933_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07806_ (.A1(\u_cpu.rf_ram.memory[48][4] ),
    .A2(_03218_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07807_ (.A1(_03222_),
    .A2(_03212_),
    .B(_03223_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07808_ (.I(_02939_),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07809_ (.A1(\u_cpu.rf_ram.memory[48][5] ),
    .A2(_03218_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07810_ (.A1(_03224_),
    .A2(_03213_),
    .B(_03225_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07811_ (.I(_02945_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07812_ (.A1(\u_cpu.rf_ram.memory[48][6] ),
    .A2(_03218_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07813_ (.A1(_03226_),
    .A2(_03213_),
    .B(_03227_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07814_ (.I(_02951_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07815_ (.A1(\u_cpu.rf_ram.memory[48][7] ),
    .A2(_03211_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07816_ (.A1(_03228_),
    .A2(_03213_),
    .B(_03229_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07817_ (.A1(_03051_),
    .A2(_03081_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07818_ (.I(_03230_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07819_ (.A1(_03181_),
    .A2(_03231_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07820_ (.I(_03232_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07821_ (.I(_03232_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07822_ (.A1(\u_cpu.rf_ram.memory[47][0] ),
    .A2(_03234_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07823_ (.A1(_03210_),
    .A2(_03233_),
    .B(_03235_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07824_ (.A1(\u_cpu.rf_ram.memory[47][1] ),
    .A2(_03234_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07825_ (.A1(_03215_),
    .A2(_03233_),
    .B(_03236_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07826_ (.I(_03232_),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07827_ (.A1(\u_cpu.rf_ram.memory[47][2] ),
    .A2(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07828_ (.A1(_03217_),
    .A2(_03233_),
    .B(_03238_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07829_ (.A1(\u_cpu.rf_ram.memory[47][3] ),
    .A2(_03237_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07830_ (.A1(_03220_),
    .A2(_03233_),
    .B(_03239_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07831_ (.A1(\u_cpu.rf_ram.memory[47][4] ),
    .A2(_03237_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07832_ (.A1(_03222_),
    .A2(_03233_),
    .B(_03240_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07833_ (.A1(\u_cpu.rf_ram.memory[47][5] ),
    .A2(_03237_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07834_ (.A1(_03224_),
    .A2(_03234_),
    .B(_03241_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07835_ (.A1(\u_cpu.rf_ram.memory[47][6] ),
    .A2(_03237_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07836_ (.A1(_03226_),
    .A2(_03234_),
    .B(_03242_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07837_ (.A1(\u_cpu.rf_ram.memory[47][7] ),
    .A2(_03232_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07838_ (.A1(_03228_),
    .A2(_03234_),
    .B(_03243_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07839_ (.A1(_02891_),
    .A2(_03168_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07840_ (.I(_03244_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07841_ (.I(_03244_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07842_ (.A1(\u_cpu.rf_ram.memory[50][0] ),
    .A2(_03246_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07843_ (.A1(_03210_),
    .A2(_03245_),
    .B(_03247_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07844_ (.A1(\u_cpu.rf_ram.memory[50][1] ),
    .A2(_03246_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07845_ (.A1(_03215_),
    .A2(_03245_),
    .B(_03248_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07846_ (.I(_03244_),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07847_ (.A1(\u_cpu.rf_ram.memory[50][2] ),
    .A2(_03249_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07848_ (.A1(_03217_),
    .A2(_03245_),
    .B(_03250_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07849_ (.A1(\u_cpu.rf_ram.memory[50][3] ),
    .A2(_03249_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07850_ (.A1(_03220_),
    .A2(_03245_),
    .B(_03251_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07851_ (.A1(\u_cpu.rf_ram.memory[50][4] ),
    .A2(_03249_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07852_ (.A1(_03222_),
    .A2(_03245_),
    .B(_03252_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07853_ (.A1(\u_cpu.rf_ram.memory[50][5] ),
    .A2(_03249_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07854_ (.A1(_03224_),
    .A2(_03246_),
    .B(_03253_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07855_ (.A1(\u_cpu.rf_ram.memory[50][6] ),
    .A2(_03249_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07856_ (.A1(_03226_),
    .A2(_03246_),
    .B(_03254_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07857_ (.A1(\u_cpu.rf_ram.memory[50][7] ),
    .A2(_03244_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07858_ (.A1(_03228_),
    .A2(_03246_),
    .B(_03255_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07859_ (.I(_03036_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07860_ (.A1(_03013_),
    .A2(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07861_ (.I(_03257_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07862_ (.I(_03258_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07863_ (.I(_03258_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07864_ (.A1(\u_cpu.rf_ram.memory[4][0] ),
    .A2(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07865_ (.A1(_02908_),
    .A2(_03259_),
    .B(_03261_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07866_ (.A1(\u_cpu.rf_ram.memory[4][1] ),
    .A2(_03260_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07867_ (.A1(_02915_),
    .A2(_03259_),
    .B(_03262_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07868_ (.I(_03258_),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07869_ (.A1(\u_cpu.rf_ram.memory[4][2] ),
    .A2(_03263_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07870_ (.A1(_02921_),
    .A2(_03259_),
    .B(_03264_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07871_ (.A1(\u_cpu.rf_ram.memory[4][3] ),
    .A2(_03263_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07872_ (.A1(_02928_),
    .A2(_03259_),
    .B(_03265_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07873_ (.A1(\u_cpu.rf_ram.memory[4][4] ),
    .A2(_03263_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07874_ (.A1(_02934_),
    .A2(_03259_),
    .B(_03266_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07875_ (.A1(\u_cpu.rf_ram.memory[4][5] ),
    .A2(_03263_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07876_ (.A1(_02940_),
    .A2(_03260_),
    .B(_03267_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07877_ (.A1(\u_cpu.rf_ram.memory[4][6] ),
    .A2(_03263_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07878_ (.A1(_02946_),
    .A2(_03260_),
    .B(_03268_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07879_ (.A1(\u_cpu.rf_ram.memory[4][7] ),
    .A2(_03258_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07880_ (.A1(_02952_),
    .A2(_03260_),
    .B(_03269_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07881_ (.I(net2),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07882_ (.I(_03270_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07883_ (.I(_03271_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07884_ (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07885_ (.I(_02726_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07886_ (.I(_03274_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07887_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_02702_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07888_ (.A1(_03275_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .B(_03276_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07889_ (.I(_03277_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07890_ (.A1(_03273_),
    .A2(\u_cpu.cpu.state.stage_two_req ),
    .B(_03278_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07891_ (.A1(_03272_),
    .A2(_03279_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07892_ (.A1(_02524_),
    .A2(_02491_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07893_ (.A1(_02519_),
    .A2(_02525_),
    .Z(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07894_ (.A1(_03280_),
    .A2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _07895_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A4(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07896_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_03283_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07897_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_03284_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07898_ (.A1(_03282_),
    .A2(_03285_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07899_ (.A1(_02505_),
    .A2(_02864_),
    .B(_02528_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07900_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07901_ (.A1(_03286_),
    .A2(_03288_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07902_ (.A1(_02495_),
    .A2(_02522_),
    .A3(_03289_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07903_ (.A1(_02632_),
    .A2(_02623_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07904_ (.A1(_02557_),
    .A2(_03290_),
    .B(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07905_ (.A1(_03273_),
    .A2(_02619_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07906_ (.A1(_02616_),
    .A2(_03292_),
    .B(_03293_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07907_ (.A1(_03279_),
    .A2(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07908_ (.A1(_02885_),
    .A2(_03295_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07909_ (.A1(_02885_),
    .A2(\u_cpu.rf_ram_if.rcnt[2] ),
    .A3(\u_cpu.rf_ram_if.rcnt[1] ),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07910_ (.A1(_02886_),
    .A2(_03295_),
    .A3(_03296_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07911_ (.A1(_01753_),
    .A2(_03296_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07912_ (.A1(_01753_),
    .A2(_03296_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07913_ (.A1(_03279_),
    .A2(_03294_),
    .A3(_03297_),
    .A4(_03298_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07914_ (.I(_03299_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07915_ (.A1(_01754_),
    .A2(_03297_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07916_ (.A1(_03295_),
    .A2(_03300_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07917_ (.A1(_02964_),
    .A2(_03068_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07918_ (.I(_03301_),
    .Z(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07919_ (.I(_03301_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07920_ (.A1(\u_cpu.rf_ram.memory[16][0] ),
    .A2(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07921_ (.A1(_03210_),
    .A2(_03302_),
    .B(_03304_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07922_ (.A1(\u_cpu.rf_ram.memory[16][1] ),
    .A2(_03303_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07923_ (.A1(_03215_),
    .A2(_03302_),
    .B(_03305_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07924_ (.I(_03301_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07925_ (.A1(\u_cpu.rf_ram.memory[16][2] ),
    .A2(_03306_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07926_ (.A1(_03217_),
    .A2(_03302_),
    .B(_03307_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07927_ (.A1(\u_cpu.rf_ram.memory[16][3] ),
    .A2(_03306_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07928_ (.A1(_03220_),
    .A2(_03302_),
    .B(_03308_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07929_ (.A1(\u_cpu.rf_ram.memory[16][4] ),
    .A2(_03306_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07930_ (.A1(_03222_),
    .A2(_03302_),
    .B(_03309_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07931_ (.A1(\u_cpu.rf_ram.memory[16][5] ),
    .A2(_03306_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07932_ (.A1(_03224_),
    .A2(_03303_),
    .B(_03310_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07933_ (.A1(\u_cpu.rf_ram.memory[16][6] ),
    .A2(_03306_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07934_ (.A1(_03226_),
    .A2(_03303_),
    .B(_03311_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07935_ (.A1(\u_cpu.rf_ram.memory[16][7] ),
    .A2(_03301_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07936_ (.A1(_03228_),
    .A2(_03303_),
    .B(_03312_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07937_ (.A1(_02964_),
    .A2(_02985_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07938_ (.I(_03313_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07939_ (.I(_03313_),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07940_ (.A1(\u_cpu.rf_ram.memory[17][0] ),
    .A2(_03315_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07941_ (.A1(_03210_),
    .A2(_03314_),
    .B(_03316_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07942_ (.A1(\u_cpu.rf_ram.memory[17][1] ),
    .A2(_03315_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07943_ (.A1(_03215_),
    .A2(_03314_),
    .B(_03317_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07944_ (.I(_03313_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07945_ (.A1(\u_cpu.rf_ram.memory[17][2] ),
    .A2(_03318_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07946_ (.A1(_03217_),
    .A2(_03314_),
    .B(_03319_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07947_ (.A1(\u_cpu.rf_ram.memory[17][3] ),
    .A2(_03318_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07948_ (.A1(_03220_),
    .A2(_03314_),
    .B(_03320_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07949_ (.A1(\u_cpu.rf_ram.memory[17][4] ),
    .A2(_03318_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07950_ (.A1(_03222_),
    .A2(_03314_),
    .B(_03321_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07951_ (.A1(\u_cpu.rf_ram.memory[17][5] ),
    .A2(_03318_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07952_ (.A1(_03224_),
    .A2(_03315_),
    .B(_03322_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07953_ (.A1(\u_cpu.rf_ram.memory[17][6] ),
    .A2(_03318_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07954_ (.A1(_03226_),
    .A2(_03315_),
    .B(_03323_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07955_ (.A1(\u_cpu.rf_ram.memory[17][7] ),
    .A2(_03313_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07956_ (.A1(_03228_),
    .A2(_03315_),
    .B(_03324_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07957_ (.I(_02906_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07958_ (.I(_03325_),
    .Z(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07959_ (.A1(_03011_),
    .A2(_03100_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07960_ (.I(_03327_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07961_ (.A1(_03181_),
    .A2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07962_ (.I(_03329_),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07963_ (.I(_03329_),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07964_ (.A1(\u_cpu.rf_ram.memory[40][0] ),
    .A2(_03331_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07965_ (.A1(_03326_),
    .A2(_03330_),
    .B(_03332_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07966_ (.I(_02913_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07967_ (.I(_03333_),
    .Z(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07968_ (.A1(\u_cpu.rf_ram.memory[40][1] ),
    .A2(_03331_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07969_ (.A1(_03334_),
    .A2(_03330_),
    .B(_03335_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07970_ (.I(_02919_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07971_ (.I(_03336_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07972_ (.I(_03329_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07973_ (.A1(\u_cpu.rf_ram.memory[40][2] ),
    .A2(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07974_ (.A1(_03337_),
    .A2(_03330_),
    .B(_03339_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07975_ (.I(_02926_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07976_ (.I(_03340_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(\u_cpu.rf_ram.memory[40][3] ),
    .A2(_03338_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07978_ (.A1(_03341_),
    .A2(_03330_),
    .B(_03342_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07979_ (.I(_02932_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07980_ (.I(_03343_),
    .Z(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07981_ (.A1(\u_cpu.rf_ram.memory[40][4] ),
    .A2(_03338_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07982_ (.A1(_03344_),
    .A2(_03330_),
    .B(_03345_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07983_ (.I(_02938_),
    .Z(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07984_ (.I(_03346_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07985_ (.A1(\u_cpu.rf_ram.memory[40][5] ),
    .A2(_03338_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07986_ (.A1(_03347_),
    .A2(_03331_),
    .B(_03348_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07987_ (.I(_02944_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07988_ (.I(_03349_),
    .Z(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07989_ (.A1(\u_cpu.rf_ram.memory[40][6] ),
    .A2(_03338_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07990_ (.A1(_03350_),
    .A2(_03331_),
    .B(_03351_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07991_ (.I(_02950_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07992_ (.I(_03352_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07993_ (.A1(\u_cpu.rf_ram.memory[40][7] ),
    .A2(_03329_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07994_ (.A1(_03353_),
    .A2(_03331_),
    .B(_03354_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07995_ (.A1(_03084_),
    .A2(_02897_),
    .A3(_03085_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07996_ (.I(_03355_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07997_ (.A1(_03053_),
    .A2(_03356_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07998_ (.I(_03357_),
    .Z(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07999_ (.I(_03357_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08000_ (.A1(\u_cpu.rf_ram.memory[119][0] ),
    .A2(_03359_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08001_ (.A1(_03326_),
    .A2(_03358_),
    .B(_03360_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08002_ (.A1(\u_cpu.rf_ram.memory[119][1] ),
    .A2(_03359_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08003_ (.A1(_03334_),
    .A2(_03358_),
    .B(_03361_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08004_ (.I(_03357_),
    .Z(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08005_ (.A1(\u_cpu.rf_ram.memory[119][2] ),
    .A2(_03362_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08006_ (.A1(_03337_),
    .A2(_03358_),
    .B(_03363_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08007_ (.A1(\u_cpu.rf_ram.memory[119][3] ),
    .A2(_03362_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08008_ (.A1(_03341_),
    .A2(_03358_),
    .B(_03364_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08009_ (.A1(\u_cpu.rf_ram.memory[119][4] ),
    .A2(_03362_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08010_ (.A1(_03344_),
    .A2(_03358_),
    .B(_03365_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08011_ (.A1(\u_cpu.rf_ram.memory[119][5] ),
    .A2(_03362_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08012_ (.A1(_03347_),
    .A2(_03359_),
    .B(_03366_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08013_ (.A1(\u_cpu.rf_ram.memory[119][6] ),
    .A2(_03362_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08014_ (.A1(_03350_),
    .A2(_03359_),
    .B(_03367_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08015_ (.A1(\u_cpu.rf_ram.memory[119][7] ),
    .A2(_03357_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08016_ (.A1(_03353_),
    .A2(_03359_),
    .B(_03368_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08017_ (.A1(_02892_),
    .A2(_02962_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08018_ (.I(_03369_),
    .Z(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08019_ (.A1(_02985_),
    .A2(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08020_ (.I(_03371_),
    .Z(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08021_ (.I(_03371_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08022_ (.A1(\u_cpu.rf_ram.memory[129][0] ),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08023_ (.A1(_03326_),
    .A2(_03372_),
    .B(_03374_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08024_ (.A1(\u_cpu.rf_ram.memory[129][1] ),
    .A2(_03373_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08025_ (.A1(_03334_),
    .A2(_03372_),
    .B(_03375_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08026_ (.I(_03371_),
    .Z(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08027_ (.A1(\u_cpu.rf_ram.memory[129][2] ),
    .A2(_03376_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08028_ (.A1(_03337_),
    .A2(_03372_),
    .B(_03377_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08029_ (.A1(\u_cpu.rf_ram.memory[129][3] ),
    .A2(_03376_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08030_ (.A1(_03341_),
    .A2(_03372_),
    .B(_03378_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08031_ (.A1(\u_cpu.rf_ram.memory[129][4] ),
    .A2(_03376_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08032_ (.A1(_03344_),
    .A2(_03372_),
    .B(_03379_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08033_ (.A1(\u_cpu.rf_ram.memory[129][5] ),
    .A2(_03376_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08034_ (.A1(_03347_),
    .A2(_03373_),
    .B(_03380_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08035_ (.A1(\u_cpu.rf_ram.memory[129][6] ),
    .A2(_03376_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08036_ (.A1(_03350_),
    .A2(_03373_),
    .B(_03381_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08037_ (.A1(\u_cpu.rf_ram.memory[129][7] ),
    .A2(_03371_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08038_ (.A1(_03353_),
    .A2(_03373_),
    .B(_03382_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08039_ (.A1(_03196_),
    .A2(_03370_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08040_ (.I(_03383_),
    .Z(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08041_ (.I(_03383_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08042_ (.A1(\u_cpu.rf_ram.memory[139][0] ),
    .A2(_03385_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08043_ (.A1(_03326_),
    .A2(_03384_),
    .B(_03386_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08044_ (.A1(\u_cpu.rf_ram.memory[139][1] ),
    .A2(_03385_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08045_ (.A1(_03334_),
    .A2(_03384_),
    .B(_03387_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08046_ (.I(_03383_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08047_ (.A1(\u_cpu.rf_ram.memory[139][2] ),
    .A2(_03388_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08048_ (.A1(_03337_),
    .A2(_03384_),
    .B(_03389_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08049_ (.A1(\u_cpu.rf_ram.memory[139][3] ),
    .A2(_03388_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08050_ (.A1(_03341_),
    .A2(_03384_),
    .B(_03390_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08051_ (.A1(\u_cpu.rf_ram.memory[139][4] ),
    .A2(_03388_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08052_ (.A1(_03344_),
    .A2(_03384_),
    .B(_03391_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08053_ (.A1(\u_cpu.rf_ram.memory[139][5] ),
    .A2(_03388_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08054_ (.A1(_03347_),
    .A2(_03385_),
    .B(_03392_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08055_ (.A1(\u_cpu.rf_ram.memory[139][6] ),
    .A2(_03388_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08056_ (.A1(_03350_),
    .A2(_03385_),
    .B(_03393_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08057_ (.A1(\u_cpu.rf_ram.memory[139][7] ),
    .A2(_03383_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08058_ (.A1(_03353_),
    .A2(_03385_),
    .B(_03394_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08059_ (.I(_03086_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08060_ (.A1(_03395_),
    .A2(_03132_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08061_ (.I(_03396_),
    .Z(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08062_ (.I(_03396_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(\u_cpu.rf_ram.memory[77][0] ),
    .A2(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08064_ (.A1(_03326_),
    .A2(_03397_),
    .B(_03399_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08065_ (.A1(\u_cpu.rf_ram.memory[77][1] ),
    .A2(_03398_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08066_ (.A1(_03334_),
    .A2(_03397_),
    .B(_03400_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08067_ (.I(_03396_),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08068_ (.A1(\u_cpu.rf_ram.memory[77][2] ),
    .A2(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08069_ (.A1(_03337_),
    .A2(_03397_),
    .B(_03402_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08070_ (.A1(\u_cpu.rf_ram.memory[77][3] ),
    .A2(_03401_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08071_ (.A1(_03341_),
    .A2(_03397_),
    .B(_03403_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08072_ (.A1(\u_cpu.rf_ram.memory[77][4] ),
    .A2(_03401_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08073_ (.A1(_03344_),
    .A2(_03397_),
    .B(_03404_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08074_ (.A1(\u_cpu.rf_ram.memory[77][5] ),
    .A2(_03401_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08075_ (.A1(_03347_),
    .A2(_03398_),
    .B(_03405_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08076_ (.A1(\u_cpu.rf_ram.memory[77][6] ),
    .A2(_03401_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08077_ (.A1(_03350_),
    .A2(_03398_),
    .B(_03406_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08078_ (.A1(\u_cpu.rf_ram.memory[77][7] ),
    .A2(_03396_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08079_ (.A1(_03353_),
    .A2(_03398_),
    .B(_03407_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08080_ (.I(_03325_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08081_ (.A1(_03395_),
    .A2(_03102_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08082_ (.I(_03409_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08083_ (.I(_03409_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08084_ (.A1(\u_cpu.rf_ram.memory[74][0] ),
    .A2(_03411_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08085_ (.A1(_03408_),
    .A2(_03410_),
    .B(_03412_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08086_ (.I(_03333_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08087_ (.A1(\u_cpu.rf_ram.memory[74][1] ),
    .A2(_03411_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08088_ (.A1(_03413_),
    .A2(_03410_),
    .B(_03414_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08089_ (.I(_03336_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08090_ (.I(_03409_),
    .Z(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08091_ (.A1(\u_cpu.rf_ram.memory[74][2] ),
    .A2(_03416_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08092_ (.A1(_03415_),
    .A2(_03410_),
    .B(_03417_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08093_ (.I(_03340_),
    .Z(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08094_ (.A1(\u_cpu.rf_ram.memory[74][3] ),
    .A2(_03416_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08095_ (.A1(_03418_),
    .A2(_03410_),
    .B(_03419_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08096_ (.I(_03343_),
    .Z(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08097_ (.A1(\u_cpu.rf_ram.memory[74][4] ),
    .A2(_03416_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08098_ (.A1(_03420_),
    .A2(_03410_),
    .B(_03421_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08099_ (.I(_03346_),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(\u_cpu.rf_ram.memory[74][5] ),
    .A2(_03416_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08101_ (.A1(_03422_),
    .A2(_03411_),
    .B(_03423_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08102_ (.I(_03349_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(\u_cpu.rf_ram.memory[74][6] ),
    .A2(_03416_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08104_ (.A1(_03424_),
    .A2(_03411_),
    .B(_03425_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08105_ (.I(_03352_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08106_ (.A1(\u_cpu.rf_ram.memory[74][7] ),
    .A2(_03409_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08107_ (.A1(_03426_),
    .A2(_03411_),
    .B(_03427_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08108_ (.A1(_03395_),
    .A2(_03153_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08109_ (.I(_03428_),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08110_ (.I(_03428_),
    .Z(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08111_ (.A1(\u_cpu.rf_ram.memory[76][0] ),
    .A2(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08112_ (.A1(_03408_),
    .A2(_03429_),
    .B(_03431_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08113_ (.A1(\u_cpu.rf_ram.memory[76][1] ),
    .A2(_03430_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08114_ (.A1(_03413_),
    .A2(_03429_),
    .B(_03432_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08115_ (.I(_03428_),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08116_ (.A1(\u_cpu.rf_ram.memory[76][2] ),
    .A2(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08117_ (.A1(_03415_),
    .A2(_03429_),
    .B(_03434_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08118_ (.A1(\u_cpu.rf_ram.memory[76][3] ),
    .A2(_03433_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08119_ (.A1(_03418_),
    .A2(_03429_),
    .B(_03435_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08120_ (.A1(\u_cpu.rf_ram.memory[76][4] ),
    .A2(_03433_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08121_ (.A1(_03420_),
    .A2(_03429_),
    .B(_03436_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08122_ (.A1(\u_cpu.rf_ram.memory[76][5] ),
    .A2(_03433_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08123_ (.A1(_03422_),
    .A2(_03430_),
    .B(_03437_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08124_ (.A1(\u_cpu.rf_ram.memory[76][6] ),
    .A2(_03433_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08125_ (.A1(_03424_),
    .A2(_03430_),
    .B(_03438_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08126_ (.A1(\u_cpu.rf_ram.memory[76][7] ),
    .A2(_03428_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08127_ (.A1(_03426_),
    .A2(_03430_),
    .B(_03439_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08128_ (.I(_03086_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08129_ (.A1(_03440_),
    .A2(_03197_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08130_ (.I(_03441_),
    .Z(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08131_ (.I(_03441_),
    .Z(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08132_ (.A1(\u_cpu.rf_ram.memory[75][0] ),
    .A2(_03443_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08133_ (.A1(_03408_),
    .A2(_03442_),
    .B(_03444_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08134_ (.A1(\u_cpu.rf_ram.memory[75][1] ),
    .A2(_03443_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08135_ (.A1(_03413_),
    .A2(_03442_),
    .B(_03445_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08136_ (.I(_03441_),
    .Z(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08137_ (.A1(\u_cpu.rf_ram.memory[75][2] ),
    .A2(_03446_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08138_ (.A1(_03415_),
    .A2(_03442_),
    .B(_03447_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08139_ (.A1(\u_cpu.rf_ram.memory[75][3] ),
    .A2(_03446_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08140_ (.A1(_03418_),
    .A2(_03442_),
    .B(_03448_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08141_ (.A1(\u_cpu.rf_ram.memory[75][4] ),
    .A2(_03446_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08142_ (.A1(_03420_),
    .A2(_03442_),
    .B(_03449_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08143_ (.A1(\u_cpu.rf_ram.memory[75][5] ),
    .A2(_03446_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08144_ (.A1(_03422_),
    .A2(_03443_),
    .B(_03450_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08145_ (.A1(\u_cpu.rf_ram.memory[75][6] ),
    .A2(_03446_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08146_ (.A1(_03424_),
    .A2(_03443_),
    .B(_03451_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08147_ (.A1(\u_cpu.rf_ram.memory[75][7] ),
    .A2(_03441_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08148_ (.A1(_03426_),
    .A2(_03443_),
    .B(_03452_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08149_ (.A1(_02889_),
    .A2(_02959_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08150_ (.I(_03453_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08151_ (.A1(_03050_),
    .A2(_03454_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08152_ (.I(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08153_ (.I(_03456_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08154_ (.I(_03456_),
    .Z(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08155_ (.A1(\u_cpu.rf_ram.memory[6][0] ),
    .A2(_03458_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08156_ (.A1(_02908_),
    .A2(_03457_),
    .B(_03459_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08157_ (.A1(\u_cpu.rf_ram.memory[6][1] ),
    .A2(_03458_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08158_ (.A1(_02915_),
    .A2(_03457_),
    .B(_03460_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08159_ (.I(_03456_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08160_ (.A1(\u_cpu.rf_ram.memory[6][2] ),
    .A2(_03461_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08161_ (.A1(_02921_),
    .A2(_03457_),
    .B(_03462_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08162_ (.A1(\u_cpu.rf_ram.memory[6][3] ),
    .A2(_03461_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08163_ (.A1(_02928_),
    .A2(_03457_),
    .B(_03463_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08164_ (.A1(\u_cpu.rf_ram.memory[6][4] ),
    .A2(_03461_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08165_ (.A1(_02934_),
    .A2(_03457_),
    .B(_03464_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08166_ (.A1(\u_cpu.rf_ram.memory[6][5] ),
    .A2(_03461_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08167_ (.A1(_02940_),
    .A2(_03458_),
    .B(_03465_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08168_ (.A1(\u_cpu.rf_ram.memory[6][6] ),
    .A2(_03461_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08169_ (.A1(_02946_),
    .A2(_03458_),
    .B(_03466_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08170_ (.A1(\u_cpu.rf_ram.memory[6][7] ),
    .A2(_03456_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08171_ (.A1(_02952_),
    .A2(_03458_),
    .B(_03467_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08172_ (.A1(_03013_),
    .A2(_03087_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08173_ (.I(_03468_),
    .Z(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08174_ (.I(_03468_),
    .Z(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08175_ (.A1(\u_cpu.rf_ram.memory[68][0] ),
    .A2(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08176_ (.A1(_03408_),
    .A2(_03469_),
    .B(_03471_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08177_ (.A1(\u_cpu.rf_ram.memory[68][1] ),
    .A2(_03470_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08178_ (.A1(_03413_),
    .A2(_03469_),
    .B(_03472_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08179_ (.I(_03468_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08180_ (.A1(\u_cpu.rf_ram.memory[68][2] ),
    .A2(_03473_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08181_ (.A1(_03415_),
    .A2(_03469_),
    .B(_03474_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08182_ (.A1(\u_cpu.rf_ram.memory[68][3] ),
    .A2(_03473_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08183_ (.A1(_03418_),
    .A2(_03469_),
    .B(_03475_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08184_ (.A1(\u_cpu.rf_ram.memory[68][4] ),
    .A2(_03473_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08185_ (.A1(_03420_),
    .A2(_03469_),
    .B(_03476_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08186_ (.A1(\u_cpu.rf_ram.memory[68][5] ),
    .A2(_03473_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08187_ (.A1(_03422_),
    .A2(_03470_),
    .B(_03477_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08188_ (.A1(\u_cpu.rf_ram.memory[68][6] ),
    .A2(_03473_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08189_ (.A1(_03424_),
    .A2(_03470_),
    .B(_03478_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08190_ (.A1(\u_cpu.rf_ram.memory[68][7] ),
    .A2(_03468_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08191_ (.A1(_03426_),
    .A2(_03470_),
    .B(_03479_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08192_ (.I(_03166_),
    .Z(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08193_ (.A1(_03440_),
    .A2(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08194_ (.I(_03481_),
    .Z(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08195_ (.I(_03481_),
    .Z(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08196_ (.A1(\u_cpu.rf_ram.memory[67][0] ),
    .A2(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08197_ (.A1(_03408_),
    .A2(_03482_),
    .B(_03484_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08198_ (.A1(\u_cpu.rf_ram.memory[67][1] ),
    .A2(_03483_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08199_ (.A1(_03413_),
    .A2(_03482_),
    .B(_03485_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08200_ (.I(_03481_),
    .Z(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08201_ (.A1(\u_cpu.rf_ram.memory[67][2] ),
    .A2(_03486_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08202_ (.A1(_03415_),
    .A2(_03482_),
    .B(_03487_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08203_ (.A1(\u_cpu.rf_ram.memory[67][3] ),
    .A2(_03486_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08204_ (.A1(_03418_),
    .A2(_03482_),
    .B(_03488_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08205_ (.A1(\u_cpu.rf_ram.memory[67][4] ),
    .A2(_03486_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08206_ (.A1(_03420_),
    .A2(_03482_),
    .B(_03489_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08207_ (.A1(\u_cpu.rf_ram.memory[67][5] ),
    .A2(_03486_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08208_ (.A1(_03422_),
    .A2(_03483_),
    .B(_03490_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08209_ (.A1(\u_cpu.rf_ram.memory[67][6] ),
    .A2(_03486_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08210_ (.A1(_03424_),
    .A2(_03483_),
    .B(_03491_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08211_ (.A1(\u_cpu.rf_ram.memory[67][7] ),
    .A2(_03481_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08212_ (.A1(_03426_),
    .A2(_03483_),
    .B(_03492_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08213_ (.I(_03325_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08214_ (.A1(_02891_),
    .A2(_03087_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08215_ (.I(_03494_),
    .Z(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08216_ (.I(_03494_),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08217_ (.A1(\u_cpu.rf_ram.memory[66][0] ),
    .A2(_03496_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08218_ (.A1(_03493_),
    .A2(_03495_),
    .B(_03497_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08219_ (.I(_03333_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08220_ (.A1(\u_cpu.rf_ram.memory[66][1] ),
    .A2(_03496_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08221_ (.A1(_03498_),
    .A2(_03495_),
    .B(_03499_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08222_ (.I(_03336_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08223_ (.I(_03494_),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08224_ (.A1(\u_cpu.rf_ram.memory[66][2] ),
    .A2(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08225_ (.A1(_03500_),
    .A2(_03495_),
    .B(_03502_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08226_ (.I(_03340_),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08227_ (.A1(\u_cpu.rf_ram.memory[66][3] ),
    .A2(_03501_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08228_ (.A1(_03503_),
    .A2(_03495_),
    .B(_03504_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08229_ (.I(_03343_),
    .Z(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08230_ (.A1(\u_cpu.rf_ram.memory[66][4] ),
    .A2(_03501_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08231_ (.A1(_03505_),
    .A2(_03495_),
    .B(_03506_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08232_ (.I(_03346_),
    .Z(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08233_ (.A1(\u_cpu.rf_ram.memory[66][5] ),
    .A2(_03501_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08234_ (.A1(_03507_),
    .A2(_03496_),
    .B(_03508_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08235_ (.I(_03349_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08236_ (.A1(\u_cpu.rf_ram.memory[66][6] ),
    .A2(_03501_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08237_ (.A1(_03509_),
    .A2(_03496_),
    .B(_03510_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08238_ (.I(_03352_),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08239_ (.A1(\u_cpu.rf_ram.memory[66][7] ),
    .A2(_03494_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08240_ (.A1(_03511_),
    .A2(_03496_),
    .B(_03512_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08241_ (.A1(_02985_),
    .A2(_03087_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08242_ (.I(_03513_),
    .Z(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08243_ (.I(_03513_),
    .Z(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08244_ (.A1(\u_cpu.rf_ram.memory[65][0] ),
    .A2(_03515_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08245_ (.A1(_03493_),
    .A2(_03514_),
    .B(_03516_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08246_ (.A1(\u_cpu.rf_ram.memory[65][1] ),
    .A2(_03515_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08247_ (.A1(_03498_),
    .A2(_03514_),
    .B(_03517_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08248_ (.I(_03513_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08249_ (.A1(\u_cpu.rf_ram.memory[65][2] ),
    .A2(_03518_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08250_ (.A1(_03500_),
    .A2(_03514_),
    .B(_03519_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08251_ (.A1(\u_cpu.rf_ram.memory[65][3] ),
    .A2(_03518_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08252_ (.A1(_03503_),
    .A2(_03514_),
    .B(_03520_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08253_ (.A1(\u_cpu.rf_ram.memory[65][4] ),
    .A2(_03518_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08254_ (.A1(_03505_),
    .A2(_03514_),
    .B(_03521_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08255_ (.A1(\u_cpu.rf_ram.memory[65][5] ),
    .A2(_03518_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08256_ (.A1(_03507_),
    .A2(_03515_),
    .B(_03522_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08257_ (.A1(\u_cpu.rf_ram.memory[65][6] ),
    .A2(_03518_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08258_ (.A1(_03509_),
    .A2(_03515_),
    .B(_03523_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08259_ (.A1(\u_cpu.rf_ram.memory[65][7] ),
    .A2(_03513_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08260_ (.A1(_03511_),
    .A2(_03515_),
    .B(_03524_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08261_ (.A1(_03068_),
    .A2(_03087_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08262_ (.I(_03525_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08263_ (.I(_03525_),
    .Z(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08264_ (.A1(\u_cpu.rf_ram.memory[64][0] ),
    .A2(_03527_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08265_ (.A1(_03493_),
    .A2(_03526_),
    .B(_03528_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08266_ (.A1(\u_cpu.rf_ram.memory[64][1] ),
    .A2(_03527_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08267_ (.A1(_03498_),
    .A2(_03526_),
    .B(_03529_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08268_ (.I(_03525_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08269_ (.A1(\u_cpu.rf_ram.memory[64][2] ),
    .A2(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08270_ (.A1(_03500_),
    .A2(_03526_),
    .B(_03531_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08271_ (.A1(\u_cpu.rf_ram.memory[64][3] ),
    .A2(_03530_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08272_ (.A1(_03503_),
    .A2(_03526_),
    .B(_03532_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08273_ (.A1(\u_cpu.rf_ram.memory[64][4] ),
    .A2(_03530_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08274_ (.A1(_03505_),
    .A2(_03526_),
    .B(_03533_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08275_ (.A1(\u_cpu.rf_ram.memory[64][5] ),
    .A2(_03530_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08276_ (.A1(_03507_),
    .A2(_03527_),
    .B(_03534_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08277_ (.A1(\u_cpu.rf_ram.memory[64][6] ),
    .A2(_03530_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08278_ (.A1(_03509_),
    .A2(_03527_),
    .B(_03535_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08279_ (.A1(\u_cpu.rf_ram.memory[64][7] ),
    .A2(_03525_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08280_ (.A1(_03511_),
    .A2(_03527_),
    .B(_03536_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08281_ (.I(_02963_),
    .Z(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08282_ (.A1(_03537_),
    .A2(_03132_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08283_ (.I(_03538_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08284_ (.I(_03538_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08285_ (.A1(\u_cpu.rf_ram.memory[29][0] ),
    .A2(_03540_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08286_ (.A1(_03493_),
    .A2(_03539_),
    .B(_03541_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08287_ (.A1(\u_cpu.rf_ram.memory[29][1] ),
    .A2(_03540_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08288_ (.A1(_03498_),
    .A2(_03539_),
    .B(_03542_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08289_ (.I(_03538_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08290_ (.A1(\u_cpu.rf_ram.memory[29][2] ),
    .A2(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08291_ (.A1(_03500_),
    .A2(_03539_),
    .B(_03544_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08292_ (.A1(\u_cpu.rf_ram.memory[29][3] ),
    .A2(_03543_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08293_ (.A1(_03503_),
    .A2(_03539_),
    .B(_03545_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08294_ (.A1(\u_cpu.rf_ram.memory[29][4] ),
    .A2(_03543_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08295_ (.A1(_03505_),
    .A2(_03539_),
    .B(_03546_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08296_ (.A1(\u_cpu.rf_ram.memory[29][5] ),
    .A2(_03543_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08297_ (.A1(_03507_),
    .A2(_03540_),
    .B(_03547_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08298_ (.A1(\u_cpu.rf_ram.memory[29][6] ),
    .A2(_03543_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08299_ (.A1(_03509_),
    .A2(_03540_),
    .B(_03548_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08300_ (.A1(\u_cpu.rf_ram.memory[29][7] ),
    .A2(_03538_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08301_ (.A1(_03511_),
    .A2(_03540_),
    .B(_03549_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08302_ (.I(_03167_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08303_ (.A1(_03550_),
    .A2(_03231_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08304_ (.I(_03551_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08305_ (.I(_03551_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08306_ (.A1(\u_cpu.rf_ram.memory[63][0] ),
    .A2(_03553_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08307_ (.A1(_03493_),
    .A2(_03552_),
    .B(_03554_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08308_ (.A1(\u_cpu.rf_ram.memory[63][1] ),
    .A2(_03553_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08309_ (.A1(_03498_),
    .A2(_03552_),
    .B(_03555_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08310_ (.I(_03551_),
    .Z(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08311_ (.A1(\u_cpu.rf_ram.memory[63][2] ),
    .A2(_03556_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08312_ (.A1(_03500_),
    .A2(_03552_),
    .B(_03557_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08313_ (.A1(\u_cpu.rf_ram.memory[63][3] ),
    .A2(_03556_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08314_ (.A1(_03503_),
    .A2(_03552_),
    .B(_03558_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08315_ (.A1(\u_cpu.rf_ram.memory[63][4] ),
    .A2(_03556_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08316_ (.A1(_03505_),
    .A2(_03552_),
    .B(_03559_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08317_ (.A1(\u_cpu.rf_ram.memory[63][5] ),
    .A2(_03556_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08318_ (.A1(_03507_),
    .A2(_03553_),
    .B(_03560_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08319_ (.A1(\u_cpu.rf_ram.memory[63][6] ),
    .A2(_03556_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08320_ (.A1(_03509_),
    .A2(_03553_),
    .B(_03561_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08321_ (.A1(\u_cpu.rf_ram.memory[63][7] ),
    .A2(_03551_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08322_ (.A1(_03511_),
    .A2(_03553_),
    .B(_03562_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08323_ (.I(_03325_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08324_ (.A1(_03082_),
    .A2(_03168_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08325_ (.I(_03564_),
    .Z(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08326_ (.I(_03564_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08327_ (.A1(\u_cpu.rf_ram.memory[62][0] ),
    .A2(_03566_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08328_ (.A1(_03563_),
    .A2(_03565_),
    .B(_03567_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08329_ (.I(_03333_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08330_ (.A1(\u_cpu.rf_ram.memory[62][1] ),
    .A2(_03566_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08331_ (.A1(_03568_),
    .A2(_03565_),
    .B(_03569_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08332_ (.I(_03336_),
    .Z(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08333_ (.I(_03564_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08334_ (.A1(\u_cpu.rf_ram.memory[62][2] ),
    .A2(_03571_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08335_ (.A1(_03570_),
    .A2(_03565_),
    .B(_03572_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08336_ (.I(_03340_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08337_ (.A1(\u_cpu.rf_ram.memory[62][3] ),
    .A2(_03571_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08338_ (.A1(_03573_),
    .A2(_03565_),
    .B(_03574_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08339_ (.I(_03343_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08340_ (.A1(\u_cpu.rf_ram.memory[62][4] ),
    .A2(_03571_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08341_ (.A1(_03575_),
    .A2(_03565_),
    .B(_03576_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08342_ (.I(_03346_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08343_ (.A1(\u_cpu.rf_ram.memory[62][5] ),
    .A2(_03571_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08344_ (.A1(_03577_),
    .A2(_03566_),
    .B(_03578_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08345_ (.I(_03349_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08346_ (.A1(\u_cpu.rf_ram.memory[62][6] ),
    .A2(_03571_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08347_ (.A1(_03579_),
    .A2(_03566_),
    .B(_03580_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08348_ (.I(_03352_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08349_ (.A1(\u_cpu.rf_ram.memory[62][7] ),
    .A2(_03564_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08350_ (.A1(_03581_),
    .A2(_03566_),
    .B(_03582_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08351_ (.A1(_03131_),
    .A2(_03168_),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08352_ (.I(_03583_),
    .Z(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08353_ (.I(_03583_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08354_ (.A1(\u_cpu.rf_ram.memory[61][0] ),
    .A2(_03585_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08355_ (.A1(_03563_),
    .A2(_03584_),
    .B(_03586_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08356_ (.A1(\u_cpu.rf_ram.memory[61][1] ),
    .A2(_03585_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08357_ (.A1(_03568_),
    .A2(_03584_),
    .B(_03587_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08358_ (.I(_03583_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08359_ (.A1(\u_cpu.rf_ram.memory[61][2] ),
    .A2(_03588_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08360_ (.A1(_03570_),
    .A2(_03584_),
    .B(_03589_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08361_ (.A1(\u_cpu.rf_ram.memory[61][3] ),
    .A2(_03588_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08362_ (.A1(_03573_),
    .A2(_03584_),
    .B(_03590_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08363_ (.A1(\u_cpu.rf_ram.memory[61][4] ),
    .A2(_03588_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08364_ (.A1(_03575_),
    .A2(_03584_),
    .B(_03591_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08365_ (.A1(\u_cpu.rf_ram.memory[61][5] ),
    .A2(_03588_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08366_ (.A1(_03577_),
    .A2(_03585_),
    .B(_03592_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08367_ (.A1(\u_cpu.rf_ram.memory[61][6] ),
    .A2(_03588_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08368_ (.A1(_03579_),
    .A2(_03585_),
    .B(_03593_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08369_ (.A1(\u_cpu.rf_ram.memory[61][7] ),
    .A2(_03583_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08370_ (.A1(_03581_),
    .A2(_03585_),
    .B(_03594_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08371_ (.I(_03167_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08372_ (.A1(_03152_),
    .A2(_03595_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08373_ (.I(_03596_),
    .Z(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08374_ (.I(_03596_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08375_ (.A1(\u_cpu.rf_ram.memory[60][0] ),
    .A2(_03598_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08376_ (.A1(_03563_),
    .A2(_03597_),
    .B(_03599_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08377_ (.A1(\u_cpu.rf_ram.memory[60][1] ),
    .A2(_03598_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08378_ (.A1(_03568_),
    .A2(_03597_),
    .B(_03600_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08379_ (.I(_03596_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08380_ (.A1(\u_cpu.rf_ram.memory[60][2] ),
    .A2(_03601_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08381_ (.A1(_03570_),
    .A2(_03597_),
    .B(_03602_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08382_ (.A1(\u_cpu.rf_ram.memory[60][3] ),
    .A2(_03601_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08383_ (.A1(_03573_),
    .A2(_03597_),
    .B(_03603_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08384_ (.A1(\u_cpu.rf_ram.memory[60][4] ),
    .A2(_03601_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08385_ (.A1(_03575_),
    .A2(_03597_),
    .B(_03604_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08386_ (.A1(\u_cpu.rf_ram.memory[60][5] ),
    .A2(_03601_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08387_ (.A1(_03577_),
    .A2(_03598_),
    .B(_03605_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08388_ (.A1(\u_cpu.rf_ram.memory[60][6] ),
    .A2(_03601_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08389_ (.A1(_03579_),
    .A2(_03598_),
    .B(_03606_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08390_ (.A1(\u_cpu.rf_ram.memory[60][7] ),
    .A2(_03596_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08391_ (.A1(_03581_),
    .A2(_03598_),
    .B(_03607_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08392_ (.A1(_03537_),
    .A2(_03480_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08393_ (.I(_03608_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08394_ (.I(_03608_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08395_ (.A1(\u_cpu.rf_ram.memory[19][0] ),
    .A2(_03610_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08396_ (.A1(_03563_),
    .A2(_03609_),
    .B(_03611_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08397_ (.A1(\u_cpu.rf_ram.memory[19][1] ),
    .A2(_03610_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08398_ (.A1(_03568_),
    .A2(_03609_),
    .B(_03612_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08399_ (.I(_03608_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08400_ (.A1(\u_cpu.rf_ram.memory[19][2] ),
    .A2(_03613_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08401_ (.A1(_03570_),
    .A2(_03609_),
    .B(_03614_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08402_ (.A1(\u_cpu.rf_ram.memory[19][3] ),
    .A2(_03613_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08403_ (.A1(_03573_),
    .A2(_03609_),
    .B(_03615_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08404_ (.A1(\u_cpu.rf_ram.memory[19][4] ),
    .A2(_03613_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08405_ (.A1(_03575_),
    .A2(_03609_),
    .B(_03616_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08406_ (.A1(\u_cpu.rf_ram.memory[19][5] ),
    .A2(_03613_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08407_ (.A1(_03577_),
    .A2(_03610_),
    .B(_03617_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08408_ (.A1(\u_cpu.rf_ram.memory[19][6] ),
    .A2(_03613_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08409_ (.A1(_03579_),
    .A2(_03610_),
    .B(_03618_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08410_ (.A1(\u_cpu.rf_ram.memory[19][7] ),
    .A2(_03608_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08411_ (.A1(_03581_),
    .A2(_03610_),
    .B(_03619_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08412_ (.I(_02906_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08413_ (.I(_03620_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08414_ (.A1(_02961_),
    .A2(_03036_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08415_ (.I(_03622_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08416_ (.I(_03623_),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08417_ (.I(_03623_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08418_ (.A1(\u_cpu.rf_ram.memory[5][0] ),
    .A2(_03625_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08419_ (.A1(_03621_),
    .A2(_03624_),
    .B(_03626_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08420_ (.I(_02913_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08421_ (.I(_03627_),
    .Z(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08422_ (.A1(\u_cpu.rf_ram.memory[5][1] ),
    .A2(_03625_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08423_ (.A1(_03628_),
    .A2(_03624_),
    .B(_03629_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08424_ (.I(_02919_),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08425_ (.I(_03630_),
    .Z(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08426_ (.I(_03623_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08427_ (.A1(\u_cpu.rf_ram.memory[5][2] ),
    .A2(_03632_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08428_ (.A1(_03631_),
    .A2(_03624_),
    .B(_03633_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08429_ (.I(_02926_),
    .Z(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08430_ (.I(_03634_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08431_ (.A1(\u_cpu.rf_ram.memory[5][3] ),
    .A2(_03632_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08432_ (.A1(_03635_),
    .A2(_03624_),
    .B(_03636_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08433_ (.I(_02932_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08434_ (.I(_03637_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08435_ (.A1(\u_cpu.rf_ram.memory[5][4] ),
    .A2(_03632_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08436_ (.A1(_03638_),
    .A2(_03624_),
    .B(_03639_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08437_ (.I(_02938_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08438_ (.I(_03640_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08439_ (.A1(\u_cpu.rf_ram.memory[5][5] ),
    .A2(_03632_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08440_ (.A1(_03641_),
    .A2(_03625_),
    .B(_03642_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08441_ (.I(_02944_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08442_ (.I(_03643_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08443_ (.A1(\u_cpu.rf_ram.memory[5][6] ),
    .A2(_03632_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08444_ (.A1(_03644_),
    .A2(_03625_),
    .B(_03645_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08445_ (.I(_02950_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08446_ (.I(_03646_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08447_ (.A1(\u_cpu.rf_ram.memory[5][7] ),
    .A2(_03623_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08448_ (.A1(_03647_),
    .A2(_03625_),
    .B(_03648_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08449_ (.A1(_03101_),
    .A2(_03595_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08450_ (.I(_03649_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08451_ (.I(_03649_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08452_ (.A1(\u_cpu.rf_ram.memory[58][0] ),
    .A2(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08453_ (.A1(_03563_),
    .A2(_03650_),
    .B(_03652_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08454_ (.A1(\u_cpu.rf_ram.memory[58][1] ),
    .A2(_03651_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08455_ (.A1(_03568_),
    .A2(_03650_),
    .B(_03653_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08456_ (.I(_03649_),
    .Z(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08457_ (.A1(\u_cpu.rf_ram.memory[58][2] ),
    .A2(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08458_ (.A1(_03570_),
    .A2(_03650_),
    .B(_03655_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08459_ (.A1(\u_cpu.rf_ram.memory[58][3] ),
    .A2(_03654_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08460_ (.A1(_03573_),
    .A2(_03650_),
    .B(_03656_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08461_ (.A1(\u_cpu.rf_ram.memory[58][4] ),
    .A2(_03654_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08462_ (.A1(_03575_),
    .A2(_03650_),
    .B(_03657_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08463_ (.A1(\u_cpu.rf_ram.memory[58][5] ),
    .A2(_03654_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08464_ (.A1(_03577_),
    .A2(_03651_),
    .B(_03658_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08465_ (.A1(\u_cpu.rf_ram.memory[58][6] ),
    .A2(_03654_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08466_ (.A1(_03579_),
    .A2(_03651_),
    .B(_03659_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08467_ (.A1(\u_cpu.rf_ram.memory[58][7] ),
    .A2(_03649_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08468_ (.A1(_03581_),
    .A2(_03651_),
    .B(_03660_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08469_ (.I(_03325_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08470_ (.A1(_03550_),
    .A2(_03183_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08471_ (.I(_03662_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08472_ (.I(_03662_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08473_ (.A1(\u_cpu.rf_ram.memory[57][0] ),
    .A2(_03664_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08474_ (.A1(_03661_),
    .A2(_03663_),
    .B(_03665_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08475_ (.I(_03333_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08476_ (.A1(\u_cpu.rf_ram.memory[57][1] ),
    .A2(_03664_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08477_ (.A1(_03666_),
    .A2(_03663_),
    .B(_03667_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08478_ (.I(_03336_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08479_ (.I(_03662_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08480_ (.A1(\u_cpu.rf_ram.memory[57][2] ),
    .A2(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08481_ (.A1(_03668_),
    .A2(_03663_),
    .B(_03670_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08482_ (.I(_03340_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08483_ (.A1(\u_cpu.rf_ram.memory[57][3] ),
    .A2(_03669_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08484_ (.A1(_03671_),
    .A2(_03663_),
    .B(_03672_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08485_ (.I(_03343_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08486_ (.A1(\u_cpu.rf_ram.memory[57][4] ),
    .A2(_03669_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08487_ (.A1(_03673_),
    .A2(_03663_),
    .B(_03674_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08488_ (.I(_03346_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08489_ (.A1(\u_cpu.rf_ram.memory[57][5] ),
    .A2(_03669_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08490_ (.A1(_03675_),
    .A2(_03664_),
    .B(_03676_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08491_ (.I(_03349_),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08492_ (.A1(\u_cpu.rf_ram.memory[57][6] ),
    .A2(_03669_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08493_ (.A1(_03677_),
    .A2(_03664_),
    .B(_03678_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08494_ (.I(_03352_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08495_ (.A1(\u_cpu.rf_ram.memory[57][7] ),
    .A2(_03662_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08496_ (.A1(_03679_),
    .A2(_03664_),
    .B(_03680_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08497_ (.A1(_03550_),
    .A2(_03328_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08498_ (.I(_03681_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08499_ (.I(_03681_),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08500_ (.A1(\u_cpu.rf_ram.memory[56][0] ),
    .A2(_03683_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08501_ (.A1(_03661_),
    .A2(_03682_),
    .B(_03684_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08502_ (.A1(\u_cpu.rf_ram.memory[56][1] ),
    .A2(_03683_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08503_ (.A1(_03666_),
    .A2(_03682_),
    .B(_03685_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08504_ (.I(_03681_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08505_ (.A1(\u_cpu.rf_ram.memory[56][2] ),
    .A2(_03686_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08506_ (.A1(_03668_),
    .A2(_03682_),
    .B(_03687_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08507_ (.A1(\u_cpu.rf_ram.memory[56][3] ),
    .A2(_03686_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08508_ (.A1(_03671_),
    .A2(_03682_),
    .B(_03688_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08509_ (.A1(\u_cpu.rf_ram.memory[56][4] ),
    .A2(_03686_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08510_ (.A1(_03673_),
    .A2(_03682_),
    .B(_03689_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08511_ (.A1(\u_cpu.rf_ram.memory[56][5] ),
    .A2(_03686_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08512_ (.A1(_03675_),
    .A2(_03683_),
    .B(_03690_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08513_ (.A1(\u_cpu.rf_ram.memory[56][6] ),
    .A2(_03686_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08514_ (.A1(_03677_),
    .A2(_03683_),
    .B(_03691_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08515_ (.A1(\u_cpu.rf_ram.memory[56][7] ),
    .A2(_03681_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08516_ (.A1(_03679_),
    .A2(_03683_),
    .B(_03692_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08517_ (.A1(_03053_),
    .A2(_03595_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08518_ (.I(_03693_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08519_ (.I(_03693_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08520_ (.A1(\u_cpu.rf_ram.memory[55][0] ),
    .A2(_03695_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08521_ (.A1(_03661_),
    .A2(_03694_),
    .B(_03696_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08522_ (.A1(\u_cpu.rf_ram.memory[55][1] ),
    .A2(_03695_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08523_ (.A1(_03666_),
    .A2(_03694_),
    .B(_03697_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08524_ (.I(_03693_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08525_ (.A1(\u_cpu.rf_ram.memory[55][2] ),
    .A2(_03698_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08526_ (.A1(_03668_),
    .A2(_03694_),
    .B(_03699_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08527_ (.A1(\u_cpu.rf_ram.memory[55][3] ),
    .A2(_03698_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08528_ (.A1(_03671_),
    .A2(_03694_),
    .B(_03700_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08529_ (.A1(\u_cpu.rf_ram.memory[55][4] ),
    .A2(_03698_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08530_ (.A1(_03673_),
    .A2(_03694_),
    .B(_03701_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08531_ (.A1(\u_cpu.rf_ram.memory[55][5] ),
    .A2(_03698_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08532_ (.A1(_03675_),
    .A2(_03695_),
    .B(_03702_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08533_ (.A1(\u_cpu.rf_ram.memory[55][6] ),
    .A2(_03698_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08534_ (.A1(_03677_),
    .A2(_03695_),
    .B(_03703_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08535_ (.A1(\u_cpu.rf_ram.memory[55][7] ),
    .A2(_03693_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08536_ (.A1(_03679_),
    .A2(_03695_),
    .B(_03704_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08537_ (.A1(_03550_),
    .A2(_03454_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08538_ (.I(_03705_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08539_ (.I(_03705_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08540_ (.A1(\u_cpu.rf_ram.memory[54][0] ),
    .A2(_03707_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08541_ (.A1(_03661_),
    .A2(_03706_),
    .B(_03708_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08542_ (.A1(\u_cpu.rf_ram.memory[54][1] ),
    .A2(_03707_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08543_ (.A1(_03666_),
    .A2(_03706_),
    .B(_03709_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08544_ (.I(_03705_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08545_ (.A1(\u_cpu.rf_ram.memory[54][2] ),
    .A2(_03710_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08546_ (.A1(_03668_),
    .A2(_03706_),
    .B(_03711_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08547_ (.A1(\u_cpu.rf_ram.memory[54][3] ),
    .A2(_03710_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08548_ (.A1(_03671_),
    .A2(_03706_),
    .B(_03712_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08549_ (.A1(\u_cpu.rf_ram.memory[54][4] ),
    .A2(_03710_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08550_ (.A1(_03673_),
    .A2(_03706_),
    .B(_03713_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08551_ (.A1(\u_cpu.rf_ram.memory[54][5] ),
    .A2(_03710_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08552_ (.A1(_03675_),
    .A2(_03707_),
    .B(_03714_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08553_ (.A1(\u_cpu.rf_ram.memory[54][6] ),
    .A2(_03710_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08554_ (.A1(_03677_),
    .A2(_03707_),
    .B(_03715_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08555_ (.A1(\u_cpu.rf_ram.memory[54][7] ),
    .A2(_03705_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08556_ (.A1(_03679_),
    .A2(_03707_),
    .B(_03716_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08557_ (.A1(_02961_),
    .A2(_03595_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08558_ (.I(_03717_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08559_ (.I(_03717_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08560_ (.A1(\u_cpu.rf_ram.memory[53][0] ),
    .A2(_03719_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08561_ (.A1(_03661_),
    .A2(_03718_),
    .B(_03720_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08562_ (.A1(\u_cpu.rf_ram.memory[53][1] ),
    .A2(_03719_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08563_ (.A1(_03666_),
    .A2(_03718_),
    .B(_03721_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08564_ (.I(_03717_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08565_ (.A1(\u_cpu.rf_ram.memory[53][2] ),
    .A2(_03722_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08566_ (.A1(_03668_),
    .A2(_03718_),
    .B(_03723_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08567_ (.A1(\u_cpu.rf_ram.memory[53][3] ),
    .A2(_03722_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08568_ (.A1(_03671_),
    .A2(_03718_),
    .B(_03724_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08569_ (.A1(\u_cpu.rf_ram.memory[53][4] ),
    .A2(_03722_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08570_ (.A1(_03673_),
    .A2(_03718_),
    .B(_03725_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08571_ (.A1(\u_cpu.rf_ram.memory[53][5] ),
    .A2(_03722_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08572_ (.A1(_03675_),
    .A2(_03719_),
    .B(_03726_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08573_ (.A1(\u_cpu.rf_ram.memory[53][6] ),
    .A2(_03722_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08574_ (.A1(_03677_),
    .A2(_03719_),
    .B(_03727_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08575_ (.A1(\u_cpu.rf_ram.memory[53][7] ),
    .A2(_03717_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08576_ (.A1(_03679_),
    .A2(_03719_),
    .B(_03728_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08577_ (.I(_02905_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08578_ (.I(_03729_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08579_ (.A1(_03013_),
    .A2(_03595_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08580_ (.I(_03731_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08581_ (.I(_03731_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08582_ (.A1(\u_cpu.rf_ram.memory[52][0] ),
    .A2(_03733_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08583_ (.A1(_03730_),
    .A2(_03732_),
    .B(_03734_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08584_ (.I(_02912_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08585_ (.I(_03735_),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08586_ (.A1(\u_cpu.rf_ram.memory[52][1] ),
    .A2(_03733_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08587_ (.A1(_03736_),
    .A2(_03732_),
    .B(_03737_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08588_ (.I(_02918_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08589_ (.I(_03738_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08590_ (.I(_03731_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08591_ (.A1(\u_cpu.rf_ram.memory[52][2] ),
    .A2(_03740_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08592_ (.A1(_03739_),
    .A2(_03732_),
    .B(_03741_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08593_ (.I(_02925_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08594_ (.I(_03742_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08595_ (.A1(\u_cpu.rf_ram.memory[52][3] ),
    .A2(_03740_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08596_ (.A1(_03743_),
    .A2(_03732_),
    .B(_03744_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08597_ (.I(_02931_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08598_ (.I(_03745_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08599_ (.A1(\u_cpu.rf_ram.memory[52][4] ),
    .A2(_03740_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08600_ (.A1(_03746_),
    .A2(_03732_),
    .B(_03747_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08601_ (.I(_02937_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08602_ (.I(_03748_),
    .Z(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08603_ (.A1(\u_cpu.rf_ram.memory[52][5] ),
    .A2(_03740_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08604_ (.A1(_03749_),
    .A2(_03733_),
    .B(_03750_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08605_ (.I(_02943_),
    .Z(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08606_ (.I(_03751_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08607_ (.A1(\u_cpu.rf_ram.memory[52][6] ),
    .A2(_03740_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08608_ (.A1(_03752_),
    .A2(_03733_),
    .B(_03753_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08609_ (.I(_02949_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08610_ (.I(_03754_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08611_ (.A1(\u_cpu.rf_ram.memory[52][7] ),
    .A2(_03731_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08612_ (.A1(_03755_),
    .A2(_03733_),
    .B(_03756_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08613_ (.A1(_03037_),
    .A2(_03183_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08614_ (.I(_03757_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08615_ (.I(_03757_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08616_ (.A1(\u_cpu.rf_ram.memory[9][0] ),
    .A2(_03759_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08617_ (.A1(_03621_),
    .A2(_03758_),
    .B(_03760_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08618_ (.A1(\u_cpu.rf_ram.memory[9][1] ),
    .A2(_03759_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08619_ (.A1(_03628_),
    .A2(_03758_),
    .B(_03761_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08620_ (.I(_03757_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08621_ (.A1(\u_cpu.rf_ram.memory[9][2] ),
    .A2(_03762_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08622_ (.A1(_03631_),
    .A2(_03758_),
    .B(_03763_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08623_ (.A1(\u_cpu.rf_ram.memory[9][3] ),
    .A2(_03762_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08624_ (.A1(_03635_),
    .A2(_03758_),
    .B(_03764_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08625_ (.A1(\u_cpu.rf_ram.memory[9][4] ),
    .A2(_03762_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08626_ (.A1(_03638_),
    .A2(_03758_),
    .B(_03765_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08627_ (.A1(\u_cpu.rf_ram.memory[9][5] ),
    .A2(_03762_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08628_ (.A1(_03641_),
    .A2(_03759_),
    .B(_03766_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08629_ (.A1(\u_cpu.rf_ram.memory[9][6] ),
    .A2(_03762_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08630_ (.A1(_03644_),
    .A2(_03759_),
    .B(_03767_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08631_ (.A1(\u_cpu.rf_ram.memory[9][7] ),
    .A2(_03757_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08632_ (.A1(_03647_),
    .A2(_03759_),
    .B(_03768_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08633_ (.A1(_03050_),
    .A2(_03231_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08634_ (.I(_03769_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08635_ (.I(_03770_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08636_ (.I(_03770_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08637_ (.A1(\u_cpu.rf_ram.memory[15][0] ),
    .A2(_03772_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08638_ (.A1(_03621_),
    .A2(_03771_),
    .B(_03773_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08639_ (.A1(\u_cpu.rf_ram.memory[15][1] ),
    .A2(_03772_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08640_ (.A1(_03628_),
    .A2(_03771_),
    .B(_03774_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08641_ (.I(_03770_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08642_ (.A1(\u_cpu.rf_ram.memory[15][2] ),
    .A2(_03775_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08643_ (.A1(_03631_),
    .A2(_03771_),
    .B(_03776_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08644_ (.A1(\u_cpu.rf_ram.memory[15][3] ),
    .A2(_03775_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08645_ (.A1(_03635_),
    .A2(_03771_),
    .B(_03777_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08646_ (.A1(\u_cpu.rf_ram.memory[15][4] ),
    .A2(_03775_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08647_ (.A1(_03638_),
    .A2(_03771_),
    .B(_03778_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08648_ (.A1(\u_cpu.rf_ram.memory[15][5] ),
    .A2(_03775_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08649_ (.A1(_03641_),
    .A2(_03772_),
    .B(_03779_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08650_ (.A1(\u_cpu.rf_ram.memory[15][6] ),
    .A2(_03775_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08651_ (.A1(_03644_),
    .A2(_03772_),
    .B(_03780_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08652_ (.A1(\u_cpu.rf_ram.memory[15][7] ),
    .A2(_03770_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08653_ (.A1(_03647_),
    .A2(_03772_),
    .B(_03781_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08654_ (.A1(_03082_),
    .A2(_03370_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08655_ (.I(_03782_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08656_ (.I(_03782_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08657_ (.A1(\u_cpu.rf_ram.memory[142][0] ),
    .A2(_03784_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08658_ (.A1(_03730_),
    .A2(_03783_),
    .B(_03785_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08659_ (.A1(\u_cpu.rf_ram.memory[142][1] ),
    .A2(_03784_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08660_ (.A1(_03736_),
    .A2(_03783_),
    .B(_03786_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08661_ (.I(_03782_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08662_ (.A1(\u_cpu.rf_ram.memory[142][2] ),
    .A2(_03787_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08663_ (.A1(_03739_),
    .A2(_03783_),
    .B(_03788_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08664_ (.A1(\u_cpu.rf_ram.memory[142][3] ),
    .A2(_03787_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08665_ (.A1(_03743_),
    .A2(_03783_),
    .B(_03789_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08666_ (.A1(\u_cpu.rf_ram.memory[142][4] ),
    .A2(_03787_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08667_ (.A1(_03746_),
    .A2(_03783_),
    .B(_03790_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08668_ (.A1(\u_cpu.rf_ram.memory[142][5] ),
    .A2(_03787_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08669_ (.A1(_03749_),
    .A2(_03784_),
    .B(_03791_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08670_ (.A1(\u_cpu.rf_ram.memory[142][6] ),
    .A2(_03787_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08671_ (.A1(_03752_),
    .A2(_03784_),
    .B(_03792_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08672_ (.A1(\u_cpu.rf_ram.memory[142][7] ),
    .A2(_03782_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08673_ (.A1(_03755_),
    .A2(_03784_),
    .B(_03793_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08674_ (.A1(_03131_),
    .A2(_03370_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08675_ (.I(_03794_),
    .Z(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08676_ (.I(_03794_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08677_ (.A1(\u_cpu.rf_ram.memory[141][0] ),
    .A2(_03796_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08678_ (.A1(_03730_),
    .A2(_03795_),
    .B(_03797_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08679_ (.A1(\u_cpu.rf_ram.memory[141][1] ),
    .A2(_03796_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08680_ (.A1(_03736_),
    .A2(_03795_),
    .B(_03798_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08681_ (.I(_03794_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08682_ (.A1(\u_cpu.rf_ram.memory[141][2] ),
    .A2(_03799_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08683_ (.A1(_03739_),
    .A2(_03795_),
    .B(_03800_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08684_ (.A1(\u_cpu.rf_ram.memory[141][3] ),
    .A2(_03799_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08685_ (.A1(_03743_),
    .A2(_03795_),
    .B(_03801_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08686_ (.A1(\u_cpu.rf_ram.memory[141][4] ),
    .A2(_03799_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08687_ (.A1(_03746_),
    .A2(_03795_),
    .B(_03802_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08688_ (.A1(\u_cpu.rf_ram.memory[141][5] ),
    .A2(_03799_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08689_ (.A1(_03749_),
    .A2(_03796_),
    .B(_03803_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08690_ (.A1(\u_cpu.rf_ram.memory[141][6] ),
    .A2(_03799_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08691_ (.A1(_03752_),
    .A2(_03796_),
    .B(_03804_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08692_ (.A1(\u_cpu.rf_ram.memory[141][7] ),
    .A2(_03794_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08693_ (.A1(_03755_),
    .A2(_03796_),
    .B(_03805_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08694_ (.A1(_03152_),
    .A2(_03370_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08695_ (.I(_03806_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08696_ (.I(_03806_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08697_ (.A1(\u_cpu.rf_ram.memory[140][0] ),
    .A2(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08698_ (.A1(_03730_),
    .A2(_03807_),
    .B(_03809_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08699_ (.A1(\u_cpu.rf_ram.memory[140][1] ),
    .A2(_03808_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08700_ (.A1(_03736_),
    .A2(_03807_),
    .B(_03810_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08701_ (.I(_03806_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08702_ (.A1(\u_cpu.rf_ram.memory[140][2] ),
    .A2(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08703_ (.A1(_03739_),
    .A2(_03807_),
    .B(_03812_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08704_ (.A1(\u_cpu.rf_ram.memory[140][3] ),
    .A2(_03811_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08705_ (.A1(_03743_),
    .A2(_03807_),
    .B(_03813_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08706_ (.A1(\u_cpu.rf_ram.memory[140][4] ),
    .A2(_03811_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08707_ (.A1(_03746_),
    .A2(_03807_),
    .B(_03814_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08708_ (.A1(\u_cpu.rf_ram.memory[140][5] ),
    .A2(_03811_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08709_ (.A1(_03749_),
    .A2(_03808_),
    .B(_03815_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08710_ (.A1(\u_cpu.rf_ram.memory[140][6] ),
    .A2(_03811_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08711_ (.A1(_03752_),
    .A2(_03808_),
    .B(_03816_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08712_ (.A1(\u_cpu.rf_ram.memory[140][7] ),
    .A2(_03806_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08713_ (.A1(_03755_),
    .A2(_03808_),
    .B(_03817_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08714_ (.A1(_03050_),
    .A2(_03132_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08715_ (.I(_03818_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08716_ (.I(_03819_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08717_ (.I(_03819_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08718_ (.A1(\u_cpu.rf_ram.memory[13][0] ),
    .A2(_03821_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08719_ (.A1(_03621_),
    .A2(_03820_),
    .B(_03822_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08720_ (.A1(\u_cpu.rf_ram.memory[13][1] ),
    .A2(_03821_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08721_ (.A1(_03628_),
    .A2(_03820_),
    .B(_03823_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08722_ (.I(_03819_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08723_ (.A1(\u_cpu.rf_ram.memory[13][2] ),
    .A2(_03824_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08724_ (.A1(_03631_),
    .A2(_03820_),
    .B(_03825_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08725_ (.A1(\u_cpu.rf_ram.memory[13][3] ),
    .A2(_03824_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08726_ (.A1(_03635_),
    .A2(_03820_),
    .B(_03826_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08727_ (.A1(\u_cpu.rf_ram.memory[13][4] ),
    .A2(_03824_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08728_ (.A1(_03638_),
    .A2(_03820_),
    .B(_03827_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08729_ (.A1(\u_cpu.rf_ram.memory[13][5] ),
    .A2(_03824_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08730_ (.A1(_03641_),
    .A2(_03821_),
    .B(_03828_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08731_ (.A1(\u_cpu.rf_ram.memory[13][6] ),
    .A2(_03824_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08732_ (.A1(_03644_),
    .A2(_03821_),
    .B(_03829_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08733_ (.A1(\u_cpu.rf_ram.memory[13][7] ),
    .A2(_03819_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08734_ (.A1(_03647_),
    .A2(_03821_),
    .B(_03830_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08735_ (.A1(_03440_),
    .A2(_03328_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08736_ (.I(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08737_ (.I(_03831_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08738_ (.A1(\u_cpu.rf_ram.memory[72][0] ),
    .A2(_03833_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08739_ (.A1(_03730_),
    .A2(_03832_),
    .B(_03834_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08740_ (.A1(\u_cpu.rf_ram.memory[72][1] ),
    .A2(_03833_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08741_ (.A1(_03736_),
    .A2(_03832_),
    .B(_03835_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08742_ (.I(_03831_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08743_ (.A1(\u_cpu.rf_ram.memory[72][2] ),
    .A2(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08744_ (.A1(_03739_),
    .A2(_03832_),
    .B(_03837_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08745_ (.A1(\u_cpu.rf_ram.memory[72][3] ),
    .A2(_03836_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08746_ (.A1(_03743_),
    .A2(_03832_),
    .B(_03838_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08747_ (.A1(\u_cpu.rf_ram.memory[72][4] ),
    .A2(_03836_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08748_ (.A1(_03746_),
    .A2(_03832_),
    .B(_03839_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08749_ (.A1(\u_cpu.rf_ram.memory[72][5] ),
    .A2(_03836_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08750_ (.A1(_03749_),
    .A2(_03833_),
    .B(_03840_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08751_ (.A1(\u_cpu.rf_ram.memory[72][6] ),
    .A2(_03836_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08752_ (.A1(_03752_),
    .A2(_03833_),
    .B(_03841_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08753_ (.A1(\u_cpu.rf_ram.memory[72][7] ),
    .A2(_03831_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08754_ (.A1(_03755_),
    .A2(_03833_),
    .B(_03842_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08755_ (.I(_03729_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08756_ (.A1(_03440_),
    .A2(_03183_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08757_ (.I(_03844_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08758_ (.I(_03844_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08759_ (.A1(\u_cpu.rf_ram.memory[73][0] ),
    .A2(_03846_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08760_ (.A1(_03843_),
    .A2(_03845_),
    .B(_03847_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08761_ (.I(_03735_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08762_ (.A1(\u_cpu.rf_ram.memory[73][1] ),
    .A2(_03846_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08763_ (.A1(_03848_),
    .A2(_03845_),
    .B(_03849_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08764_ (.I(_03738_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08765_ (.I(_03844_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08766_ (.A1(\u_cpu.rf_ram.memory[73][2] ),
    .A2(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08767_ (.A1(_03850_),
    .A2(_03845_),
    .B(_03852_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08768_ (.I(_03742_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08769_ (.A1(\u_cpu.rf_ram.memory[73][3] ),
    .A2(_03851_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08770_ (.A1(_03853_),
    .A2(_03845_),
    .B(_03854_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08771_ (.I(_03745_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08772_ (.A1(\u_cpu.rf_ram.memory[73][4] ),
    .A2(_03851_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08773_ (.A1(_03855_),
    .A2(_03845_),
    .B(_03856_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08774_ (.I(_03748_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08775_ (.A1(\u_cpu.rf_ram.memory[73][5] ),
    .A2(_03851_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08776_ (.A1(_03857_),
    .A2(_03846_),
    .B(_03858_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08777_ (.I(_03751_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08778_ (.A1(\u_cpu.rf_ram.memory[73][6] ),
    .A2(_03851_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08779_ (.A1(_03859_),
    .A2(_03846_),
    .B(_03860_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08780_ (.I(_03754_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08781_ (.A1(\u_cpu.rf_ram.memory[73][7] ),
    .A2(_03844_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08782_ (.A1(_03861_),
    .A2(_03846_),
    .B(_03862_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08783_ (.A1(_03052_),
    .A2(_03395_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08784_ (.I(_03863_),
    .Z(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08785_ (.I(_03863_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08786_ (.A1(\u_cpu.rf_ram.memory[71][0] ),
    .A2(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08787_ (.A1(_03843_),
    .A2(_03864_),
    .B(_03866_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08788_ (.A1(\u_cpu.rf_ram.memory[71][1] ),
    .A2(_03865_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08789_ (.A1(_03848_),
    .A2(_03864_),
    .B(_03867_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08790_ (.I(_03863_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08791_ (.A1(\u_cpu.rf_ram.memory[71][2] ),
    .A2(_03868_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08792_ (.A1(_03850_),
    .A2(_03864_),
    .B(_03869_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08793_ (.A1(\u_cpu.rf_ram.memory[71][3] ),
    .A2(_03868_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08794_ (.A1(_03853_),
    .A2(_03864_),
    .B(_03870_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08795_ (.A1(\u_cpu.rf_ram.memory[71][4] ),
    .A2(_03868_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08796_ (.A1(_03855_),
    .A2(_03864_),
    .B(_03871_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08797_ (.A1(\u_cpu.rf_ram.memory[71][5] ),
    .A2(_03868_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08798_ (.A1(_03857_),
    .A2(_03865_),
    .B(_03872_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08799_ (.A1(\u_cpu.rf_ram.memory[71][6] ),
    .A2(_03868_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08800_ (.A1(_03859_),
    .A2(_03865_),
    .B(_03873_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08801_ (.A1(\u_cpu.rf_ram.memory[71][7] ),
    .A2(_03863_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08802_ (.A1(_03861_),
    .A2(_03865_),
    .B(_03874_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08803_ (.A1(_03440_),
    .A2(_03454_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08804_ (.I(_03875_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08805_ (.I(_03875_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08806_ (.A1(\u_cpu.rf_ram.memory[70][0] ),
    .A2(_03877_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08807_ (.A1(_03843_),
    .A2(_03876_),
    .B(_03878_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08808_ (.A1(\u_cpu.rf_ram.memory[70][1] ),
    .A2(_03877_),
    .ZN(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08809_ (.A1(_03848_),
    .A2(_03876_),
    .B(_03879_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08810_ (.I(_03875_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08811_ (.A1(\u_cpu.rf_ram.memory[70][2] ),
    .A2(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08812_ (.A1(_03850_),
    .A2(_03876_),
    .B(_03881_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08813_ (.A1(\u_cpu.rf_ram.memory[70][3] ),
    .A2(_03880_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08814_ (.A1(_03853_),
    .A2(_03876_),
    .B(_03882_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08815_ (.A1(\u_cpu.rf_ram.memory[70][4] ),
    .A2(_03880_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08816_ (.A1(_03855_),
    .A2(_03876_),
    .B(_03883_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08817_ (.A1(\u_cpu.rf_ram.memory[70][5] ),
    .A2(_03880_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08818_ (.A1(_03857_),
    .A2(_03877_),
    .B(_03884_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08819_ (.A1(\u_cpu.rf_ram.memory[70][6] ),
    .A2(_03880_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08820_ (.A1(_03859_),
    .A2(_03877_),
    .B(_03885_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08821_ (.A1(\u_cpu.rf_ram.memory[70][7] ),
    .A2(_03875_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08822_ (.A1(_03861_),
    .A2(_03877_),
    .B(_03886_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08823_ (.I(_03369_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08824_ (.A1(_03230_),
    .A2(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08825_ (.I(_03888_),
    .Z(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08826_ (.I(_03888_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08827_ (.A1(\u_cpu.rf_ram.memory[143][0] ),
    .A2(_03890_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08828_ (.A1(_03843_),
    .A2(_03889_),
    .B(_03891_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08829_ (.A1(\u_cpu.rf_ram.memory[143][1] ),
    .A2(_03890_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08830_ (.A1(_03848_),
    .A2(_03889_),
    .B(_03892_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08831_ (.I(_03888_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08832_ (.A1(\u_cpu.rf_ram.memory[143][2] ),
    .A2(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08833_ (.A1(_03850_),
    .A2(_03889_),
    .B(_03894_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08834_ (.A1(\u_cpu.rf_ram.memory[143][3] ),
    .A2(_03893_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08835_ (.A1(_03853_),
    .A2(_03889_),
    .B(_03895_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08836_ (.A1(\u_cpu.rf_ram.memory[143][4] ),
    .A2(_03893_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08837_ (.A1(_03855_),
    .A2(_03889_),
    .B(_03896_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08838_ (.A1(\u_cpu.rf_ram.memory[143][5] ),
    .A2(_03893_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08839_ (.A1(_03857_),
    .A2(_03890_),
    .B(_03897_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08840_ (.A1(\u_cpu.rf_ram.memory[143][6] ),
    .A2(_03893_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08841_ (.A1(_03859_),
    .A2(_03890_),
    .B(_03898_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08842_ (.A1(\u_cpu.rf_ram.memory[143][7] ),
    .A2(_03888_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08843_ (.A1(_03861_),
    .A2(_03890_),
    .B(_03899_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08844_ (.A1(_03256_),
    .A2(_03083_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08845_ (.I(_03900_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08846_ (.I(_03901_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08847_ (.I(_03901_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08848_ (.A1(\u_cpu.rf_ram.memory[14][0] ),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08849_ (.A1(_03621_),
    .A2(_03902_),
    .B(_03904_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08850_ (.A1(\u_cpu.rf_ram.memory[14][1] ),
    .A2(_03903_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08851_ (.A1(_03628_),
    .A2(_03902_),
    .B(_03905_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08852_ (.I(_03901_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08853_ (.A1(\u_cpu.rf_ram.memory[14][2] ),
    .A2(_03906_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08854_ (.A1(_03631_),
    .A2(_03902_),
    .B(_03907_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08855_ (.A1(\u_cpu.rf_ram.memory[14][3] ),
    .A2(_03906_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08856_ (.A1(_03635_),
    .A2(_03902_),
    .B(_03908_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08857_ (.A1(\u_cpu.rf_ram.memory[14][4] ),
    .A2(_03906_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08858_ (.A1(_03638_),
    .A2(_03902_),
    .B(_03909_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08859_ (.A1(\u_cpu.rf_ram.memory[14][5] ),
    .A2(_03906_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08860_ (.A1(_03641_),
    .A2(_03903_),
    .B(_03910_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08861_ (.A1(\u_cpu.rf_ram.memory[14][6] ),
    .A2(_03906_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08862_ (.A1(_03644_),
    .A2(_03903_),
    .B(_03911_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08863_ (.A1(\u_cpu.rf_ram.memory[14][7] ),
    .A2(_03901_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08864_ (.A1(_03647_),
    .A2(_03903_),
    .B(_03912_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08865_ (.A1(_03101_),
    .A2(_03887_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08866_ (.I(_03913_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08867_ (.I(_03913_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08868_ (.A1(\u_cpu.rf_ram.memory[138][0] ),
    .A2(_03915_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08869_ (.A1(_03843_),
    .A2(_03914_),
    .B(_03916_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08870_ (.A1(\u_cpu.rf_ram.memory[138][1] ),
    .A2(_03915_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08871_ (.A1(_03848_),
    .A2(_03914_),
    .B(_03917_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08872_ (.I(_03913_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08873_ (.A1(\u_cpu.rf_ram.memory[138][2] ),
    .A2(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08874_ (.A1(_03850_),
    .A2(_03914_),
    .B(_03919_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08875_ (.A1(\u_cpu.rf_ram.memory[138][3] ),
    .A2(_03918_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08876_ (.A1(_03853_),
    .A2(_03914_),
    .B(_03920_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08877_ (.A1(\u_cpu.rf_ram.memory[138][4] ),
    .A2(_03918_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08878_ (.A1(_03855_),
    .A2(_03914_),
    .B(_03921_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08879_ (.A1(\u_cpu.rf_ram.memory[138][5] ),
    .A2(_03918_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08880_ (.A1(_03857_),
    .A2(_03915_),
    .B(_03922_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08881_ (.A1(\u_cpu.rf_ram.memory[138][6] ),
    .A2(_03918_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08882_ (.A1(_03859_),
    .A2(_03915_),
    .B(_03923_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08883_ (.A1(\u_cpu.rf_ram.memory[138][7] ),
    .A2(_03913_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08884_ (.A1(_03861_),
    .A2(_03915_),
    .B(_03924_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08885_ (.I(_03729_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08886_ (.A1(_03052_),
    .A2(_03104_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08887_ (.I(_03926_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08888_ (.I(_03926_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08889_ (.A1(\u_cpu.rf_ram.memory[39][0] ),
    .A2(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08890_ (.A1(_03925_),
    .A2(_03927_),
    .B(_03929_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08891_ (.I(_03735_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08892_ (.A1(\u_cpu.rf_ram.memory[39][1] ),
    .A2(_03928_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08893_ (.A1(_03930_),
    .A2(_03927_),
    .B(_03931_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08894_ (.I(_03738_),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08895_ (.I(_03926_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08896_ (.A1(\u_cpu.rf_ram.memory[39][2] ),
    .A2(_03933_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08897_ (.A1(_03932_),
    .A2(_03927_),
    .B(_03934_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08898_ (.I(_03742_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08899_ (.A1(\u_cpu.rf_ram.memory[39][3] ),
    .A2(_03933_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08900_ (.A1(_03935_),
    .A2(_03927_),
    .B(_03936_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08901_ (.I(_03745_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08902_ (.A1(\u_cpu.rf_ram.memory[39][4] ),
    .A2(_03933_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08903_ (.A1(_03937_),
    .A2(_03927_),
    .B(_03938_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08904_ (.I(_03748_),
    .Z(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08905_ (.A1(\u_cpu.rf_ram.memory[39][5] ),
    .A2(_03933_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08906_ (.A1(_03939_),
    .A2(_03928_),
    .B(_03940_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08907_ (.I(_03751_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08908_ (.A1(\u_cpu.rf_ram.memory[39][6] ),
    .A2(_03933_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08909_ (.A1(_03941_),
    .A2(_03928_),
    .B(_03942_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08910_ (.I(_03754_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08911_ (.A1(\u_cpu.rf_ram.memory[39][7] ),
    .A2(_03926_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08912_ (.A1(_03943_),
    .A2(_03928_),
    .B(_03944_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08913_ (.A1(_03182_),
    .A2(_03887_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08914_ (.I(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08915_ (.I(_03945_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08916_ (.A1(\u_cpu.rf_ram.memory[137][0] ),
    .A2(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08917_ (.A1(_03925_),
    .A2(_03946_),
    .B(_03948_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(\u_cpu.rf_ram.memory[137][1] ),
    .A2(_03947_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08919_ (.A1(_03930_),
    .A2(_03946_),
    .B(_03949_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08920_ (.I(_03945_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08921_ (.A1(\u_cpu.rf_ram.memory[137][2] ),
    .A2(_03950_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08922_ (.A1(_03932_),
    .A2(_03946_),
    .B(_03951_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08923_ (.A1(\u_cpu.rf_ram.memory[137][3] ),
    .A2(_03950_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08924_ (.A1(_03935_),
    .A2(_03946_),
    .B(_03952_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08925_ (.A1(\u_cpu.rf_ram.memory[137][4] ),
    .A2(_03950_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08926_ (.A1(_03937_),
    .A2(_03946_),
    .B(_03953_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08927_ (.A1(\u_cpu.rf_ram.memory[137][5] ),
    .A2(_03950_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08928_ (.A1(_03939_),
    .A2(_03947_),
    .B(_03954_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08929_ (.A1(\u_cpu.rf_ram.memory[137][6] ),
    .A2(_03950_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08930_ (.A1(_03941_),
    .A2(_03947_),
    .B(_03955_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08931_ (.A1(\u_cpu.rf_ram.memory[137][7] ),
    .A2(_03945_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08932_ (.A1(_03943_),
    .A2(_03947_),
    .B(_03956_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08933_ (.A1(_02984_),
    .A2(_03550_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08934_ (.I(_03957_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08935_ (.I(_03957_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08936_ (.A1(\u_cpu.rf_ram.memory[49][0] ),
    .A2(_03959_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08937_ (.A1(_03925_),
    .A2(_03958_),
    .B(_03960_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08938_ (.A1(\u_cpu.rf_ram.memory[49][1] ),
    .A2(_03959_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08939_ (.A1(_03930_),
    .A2(_03958_),
    .B(_03961_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08940_ (.I(_03957_),
    .Z(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08941_ (.A1(\u_cpu.rf_ram.memory[49][2] ),
    .A2(_03962_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08942_ (.A1(_03932_),
    .A2(_03958_),
    .B(_03963_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08943_ (.A1(\u_cpu.rf_ram.memory[49][3] ),
    .A2(_03962_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08944_ (.A1(_03935_),
    .A2(_03958_),
    .B(_03964_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08945_ (.A1(\u_cpu.rf_ram.memory[49][4] ),
    .A2(_03962_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08946_ (.A1(_03937_),
    .A2(_03958_),
    .B(_03965_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08947_ (.A1(\u_cpu.rf_ram.memory[49][5] ),
    .A2(_03962_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08948_ (.A1(_03939_),
    .A2(_03959_),
    .B(_03966_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08949_ (.A1(\u_cpu.rf_ram.memory[49][6] ),
    .A2(_03962_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08950_ (.A1(_03941_),
    .A2(_03959_),
    .B(_03967_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08951_ (.A1(\u_cpu.rf_ram.memory[49][7] ),
    .A2(_03957_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08952_ (.A1(_03943_),
    .A2(_03959_),
    .B(_03968_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08953_ (.A1(_03327_),
    .A2(_03887_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08954_ (.I(_03969_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08955_ (.I(_03969_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08956_ (.A1(\u_cpu.rf_ram.memory[136][0] ),
    .A2(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08957_ (.A1(_03925_),
    .A2(_03970_),
    .B(_03972_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08958_ (.A1(\u_cpu.rf_ram.memory[136][1] ),
    .A2(_03971_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08959_ (.A1(_03930_),
    .A2(_03970_),
    .B(_03973_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08960_ (.I(_03969_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08961_ (.A1(\u_cpu.rf_ram.memory[136][2] ),
    .A2(_03974_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08962_ (.A1(_03932_),
    .A2(_03970_),
    .B(_03975_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08963_ (.A1(\u_cpu.rf_ram.memory[136][3] ),
    .A2(_03974_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08964_ (.A1(_03935_),
    .A2(_03970_),
    .B(_03976_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08965_ (.A1(\u_cpu.rf_ram.memory[136][4] ),
    .A2(_03974_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08966_ (.A1(_03937_),
    .A2(_03970_),
    .B(_03977_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08967_ (.A1(\u_cpu.rf_ram.memory[136][5] ),
    .A2(_03974_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08968_ (.A1(_03939_),
    .A2(_03971_),
    .B(_03978_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08969_ (.A1(\u_cpu.rf_ram.memory[136][6] ),
    .A2(_03974_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08970_ (.A1(_03941_),
    .A2(_03971_),
    .B(_03979_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08971_ (.A1(\u_cpu.rf_ram.memory[136][7] ),
    .A2(_03969_),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08972_ (.A1(_03943_),
    .A2(_03971_),
    .B(_03980_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08973_ (.A1(_03052_),
    .A2(_03887_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08974_ (.I(_03981_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08975_ (.I(_03981_),
    .Z(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08976_ (.A1(\u_cpu.rf_ram.memory[135][0] ),
    .A2(_03983_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08977_ (.A1(_03925_),
    .A2(_03982_),
    .B(_03984_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08978_ (.A1(\u_cpu.rf_ram.memory[135][1] ),
    .A2(_03983_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08979_ (.A1(_03930_),
    .A2(_03982_),
    .B(_03985_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08980_ (.I(_03981_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08981_ (.A1(\u_cpu.rf_ram.memory[135][2] ),
    .A2(_03986_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08982_ (.A1(_03932_),
    .A2(_03982_),
    .B(_03987_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08983_ (.A1(\u_cpu.rf_ram.memory[135][3] ),
    .A2(_03986_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08984_ (.A1(_03935_),
    .A2(_03982_),
    .B(_03988_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08985_ (.A1(\u_cpu.rf_ram.memory[135][4] ),
    .A2(_03986_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08986_ (.A1(_03937_),
    .A2(_03982_),
    .B(_03989_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08987_ (.A1(\u_cpu.rf_ram.memory[135][5] ),
    .A2(_03986_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08988_ (.A1(_03939_),
    .A2(_03983_),
    .B(_03990_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08989_ (.A1(\u_cpu.rf_ram.memory[135][6] ),
    .A2(_03986_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08990_ (.A1(_03941_),
    .A2(_03983_),
    .B(_03991_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08991_ (.A1(\u_cpu.rf_ram.memory[135][7] ),
    .A2(_03981_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08992_ (.A1(_03943_),
    .A2(_03983_),
    .B(_03992_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08993_ (.I(_03729_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08994_ (.A1(_03369_),
    .A2(_03454_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08995_ (.I(_03994_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08996_ (.I(_03994_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08997_ (.A1(\u_cpu.rf_ram.memory[134][0] ),
    .A2(_03996_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08998_ (.A1(_03993_),
    .A2(_03995_),
    .B(_03997_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08999_ (.I(_03735_),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09000_ (.A1(\u_cpu.rf_ram.memory[134][1] ),
    .A2(_03996_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09001_ (.A1(_03998_),
    .A2(_03995_),
    .B(_03999_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09002_ (.I(_03738_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09003_ (.I(_03994_),
    .Z(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09004_ (.A1(\u_cpu.rf_ram.memory[134][2] ),
    .A2(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09005_ (.A1(_04000_),
    .A2(_03995_),
    .B(_04002_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09006_ (.I(_03742_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09007_ (.A1(\u_cpu.rf_ram.memory[134][3] ),
    .A2(_04001_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09008_ (.A1(_04003_),
    .A2(_03995_),
    .B(_04004_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09009_ (.I(_03745_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09010_ (.A1(\u_cpu.rf_ram.memory[134][4] ),
    .A2(_04001_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09011_ (.A1(_04005_),
    .A2(_03995_),
    .B(_04006_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09012_ (.I(_03748_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09013_ (.A1(\u_cpu.rf_ram.memory[134][5] ),
    .A2(_04001_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09014_ (.A1(_04007_),
    .A2(_03996_),
    .B(_04008_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09015_ (.I(_03751_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09016_ (.A1(\u_cpu.rf_ram.memory[134][6] ),
    .A2(_04001_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09017_ (.A1(_04009_),
    .A2(_03996_),
    .B(_04010_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09018_ (.I(_03754_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09019_ (.A1(\u_cpu.rf_ram.memory[134][7] ),
    .A2(_03994_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09020_ (.A1(_04011_),
    .A2(_03996_),
    .B(_04012_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09021_ (.I(_03369_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09022_ (.A1(_02961_),
    .A2(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09023_ (.I(_04014_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09024_ (.I(_04014_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09025_ (.A1(\u_cpu.rf_ram.memory[133][0] ),
    .A2(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09026_ (.A1(_03993_),
    .A2(_04015_),
    .B(_04017_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09027_ (.A1(\u_cpu.rf_ram.memory[133][1] ),
    .A2(_04016_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09028_ (.A1(_03998_),
    .A2(_04015_),
    .B(_04018_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09029_ (.I(_04014_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09030_ (.A1(\u_cpu.rf_ram.memory[133][2] ),
    .A2(_04019_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09031_ (.A1(_04000_),
    .A2(_04015_),
    .B(_04020_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09032_ (.A1(\u_cpu.rf_ram.memory[133][3] ),
    .A2(_04019_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09033_ (.A1(_04003_),
    .A2(_04015_),
    .B(_04021_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09034_ (.A1(\u_cpu.rf_ram.memory[133][4] ),
    .A2(_04019_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09035_ (.A1(_04005_),
    .A2(_04015_),
    .B(_04022_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09036_ (.A1(\u_cpu.rf_ram.memory[133][5] ),
    .A2(_04019_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09037_ (.A1(_04007_),
    .A2(_04016_),
    .B(_04023_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09038_ (.A1(\u_cpu.rf_ram.memory[133][6] ),
    .A2(_04019_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09039_ (.A1(_04009_),
    .A2(_04016_),
    .B(_04024_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09040_ (.A1(\u_cpu.rf_ram.memory[133][7] ),
    .A2(_04014_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09041_ (.A1(_04011_),
    .A2(_04016_),
    .B(_04025_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09042_ (.A1(_03012_),
    .A2(_04013_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09043_ (.I(_04026_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09044_ (.I(_04026_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09045_ (.A1(\u_cpu.rf_ram.memory[132][0] ),
    .A2(_04028_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09046_ (.A1(_03993_),
    .A2(_04027_),
    .B(_04029_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09047_ (.A1(\u_cpu.rf_ram.memory[132][1] ),
    .A2(_04028_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09048_ (.A1(_03998_),
    .A2(_04027_),
    .B(_04030_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09049_ (.I(_04026_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09050_ (.A1(\u_cpu.rf_ram.memory[132][2] ),
    .A2(_04031_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09051_ (.A1(_04000_),
    .A2(_04027_),
    .B(_04032_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09052_ (.A1(\u_cpu.rf_ram.memory[132][3] ),
    .A2(_04031_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09053_ (.A1(_04003_),
    .A2(_04027_),
    .B(_04033_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09054_ (.A1(\u_cpu.rf_ram.memory[132][4] ),
    .A2(_04031_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09055_ (.A1(_04005_),
    .A2(_04027_),
    .B(_04034_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09056_ (.A1(\u_cpu.rf_ram.memory[132][5] ),
    .A2(_04031_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09057_ (.A1(_04007_),
    .A2(_04028_),
    .B(_04035_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09058_ (.A1(\u_cpu.rf_ram.memory[132][6] ),
    .A2(_04031_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09059_ (.A1(_04009_),
    .A2(_04028_),
    .B(_04036_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09060_ (.A1(\u_cpu.rf_ram.memory[132][7] ),
    .A2(_04026_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09061_ (.A1(_04011_),
    .A2(_04028_),
    .B(_04037_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09062_ (.A1(_03166_),
    .A2(_04013_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09063_ (.I(_04038_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09064_ (.I(_04038_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09065_ (.A1(\u_cpu.rf_ram.memory[131][0] ),
    .A2(_04040_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09066_ (.A1(_03993_),
    .A2(_04039_),
    .B(_04041_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09067_ (.A1(\u_cpu.rf_ram.memory[131][1] ),
    .A2(_04040_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09068_ (.A1(_03998_),
    .A2(_04039_),
    .B(_04042_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09069_ (.I(_04038_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09070_ (.A1(\u_cpu.rf_ram.memory[131][2] ),
    .A2(_04043_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09071_ (.A1(_04000_),
    .A2(_04039_),
    .B(_04044_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09072_ (.A1(\u_cpu.rf_ram.memory[131][3] ),
    .A2(_04043_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09073_ (.A1(_04003_),
    .A2(_04039_),
    .B(_04045_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09074_ (.A1(\u_cpu.rf_ram.memory[131][4] ),
    .A2(_04043_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09075_ (.A1(_04005_),
    .A2(_04039_),
    .B(_04046_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09076_ (.A1(\u_cpu.rf_ram.memory[131][5] ),
    .A2(_04043_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09077_ (.A1(_04007_),
    .A2(_04040_),
    .B(_04047_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09078_ (.A1(\u_cpu.rf_ram.memory[131][6] ),
    .A2(_04043_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09079_ (.A1(_04009_),
    .A2(_04040_),
    .B(_04048_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09080_ (.A1(\u_cpu.rf_ram.memory[131][7] ),
    .A2(_04038_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09081_ (.A1(_04011_),
    .A2(_04040_),
    .B(_04049_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09082_ (.A1(_02890_),
    .A2(_04013_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09083_ (.I(_04050_),
    .Z(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09084_ (.I(_04050_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09085_ (.A1(\u_cpu.rf_ram.memory[130][0] ),
    .A2(_04052_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09086_ (.A1(_03993_),
    .A2(_04051_),
    .B(_04053_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09087_ (.A1(\u_cpu.rf_ram.memory[130][1] ),
    .A2(_04052_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09088_ (.A1(_03998_),
    .A2(_04051_),
    .B(_04054_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09089_ (.I(_04050_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09090_ (.A1(\u_cpu.rf_ram.memory[130][2] ),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09091_ (.A1(_04000_),
    .A2(_04051_),
    .B(_04056_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09092_ (.A1(\u_cpu.rf_ram.memory[130][3] ),
    .A2(_04055_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09093_ (.A1(_04003_),
    .A2(_04051_),
    .B(_04057_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09094_ (.A1(\u_cpu.rf_ram.memory[130][4] ),
    .A2(_04055_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09095_ (.A1(_04005_),
    .A2(_04051_),
    .B(_04058_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09096_ (.A1(\u_cpu.rf_ram.memory[130][5] ),
    .A2(_04055_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09097_ (.A1(_04007_),
    .A2(_04052_),
    .B(_04059_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09098_ (.A1(\u_cpu.rf_ram.memory[130][6] ),
    .A2(_04055_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09099_ (.A1(_04009_),
    .A2(_04052_),
    .B(_04060_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09100_ (.A1(\u_cpu.rf_ram.memory[130][7] ),
    .A2(_04050_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09101_ (.A1(_04011_),
    .A2(_04052_),
    .B(_04061_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09102_ (.I(_02907_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09103_ (.A1(_03256_),
    .A2(_03153_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09104_ (.I(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09105_ (.I(_04064_),
    .Z(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09106_ (.I(_04064_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09107_ (.A1(\u_cpu.rf_ram.memory[12][0] ),
    .A2(_04066_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09108_ (.A1(_04062_),
    .A2(_04065_),
    .B(_04067_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09109_ (.I(_02914_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09110_ (.A1(\u_cpu.rf_ram.memory[12][1] ),
    .A2(_04066_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09111_ (.A1(_04068_),
    .A2(_04065_),
    .B(_04069_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09112_ (.I(_02920_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09113_ (.I(_04064_),
    .Z(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09114_ (.A1(\u_cpu.rf_ram.memory[12][2] ),
    .A2(_04071_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09115_ (.A1(_04070_),
    .A2(_04065_),
    .B(_04072_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09116_ (.I(_02927_),
    .Z(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09117_ (.A1(\u_cpu.rf_ram.memory[12][3] ),
    .A2(_04071_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09118_ (.A1(_04073_),
    .A2(_04065_),
    .B(_04074_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09119_ (.I(_02933_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09120_ (.A1(\u_cpu.rf_ram.memory[12][4] ),
    .A2(_04071_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09121_ (.A1(_04075_),
    .A2(_04065_),
    .B(_04076_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09122_ (.I(_02939_),
    .Z(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09123_ (.A1(\u_cpu.rf_ram.memory[12][5] ),
    .A2(_04071_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09124_ (.A1(_04077_),
    .A2(_04066_),
    .B(_04078_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09125_ (.I(_02945_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09126_ (.A1(\u_cpu.rf_ram.memory[12][6] ),
    .A2(_04071_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09127_ (.A1(_04079_),
    .A2(_04066_),
    .B(_04080_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09128_ (.I(_02951_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09129_ (.A1(\u_cpu.rf_ram.memory[12][7] ),
    .A2(_04064_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09130_ (.A1(_04081_),
    .A2(_04066_),
    .B(_04082_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09131_ (.I(_03729_),
    .Z(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09132_ (.A1(_03537_),
    .A2(_03454_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09133_ (.I(_04084_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09134_ (.I(_04084_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09135_ (.A1(\u_cpu.rf_ram.memory[22][0] ),
    .A2(_04086_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09136_ (.A1(_04083_),
    .A2(_04085_),
    .B(_04087_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09137_ (.I(_03735_),
    .Z(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09138_ (.A1(\u_cpu.rf_ram.memory[22][1] ),
    .A2(_04086_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09139_ (.A1(_04088_),
    .A2(_04085_),
    .B(_04089_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09140_ (.I(_03738_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09141_ (.I(_04084_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09142_ (.A1(\u_cpu.rf_ram.memory[22][2] ),
    .A2(_04091_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09143_ (.A1(_04090_),
    .A2(_04085_),
    .B(_04092_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09144_ (.I(_03742_),
    .Z(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09145_ (.A1(\u_cpu.rf_ram.memory[22][3] ),
    .A2(_04091_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09146_ (.A1(_04093_),
    .A2(_04085_),
    .B(_04094_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09147_ (.I(_03745_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09148_ (.A1(\u_cpu.rf_ram.memory[22][4] ),
    .A2(_04091_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09149_ (.A1(_04095_),
    .A2(_04085_),
    .B(_04096_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09150_ (.I(_03748_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09151_ (.A1(\u_cpu.rf_ram.memory[22][5] ),
    .A2(_04091_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09152_ (.A1(_04097_),
    .A2(_04086_),
    .B(_04098_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09153_ (.I(_03751_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09154_ (.A1(\u_cpu.rf_ram.memory[22][6] ),
    .A2(_04091_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09155_ (.A1(_04099_),
    .A2(_04086_),
    .B(_04100_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09156_ (.I(_03754_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09157_ (.A1(\u_cpu.rf_ram.memory[22][7] ),
    .A2(_04084_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09158_ (.A1(_04101_),
    .A2(_04086_),
    .B(_04102_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09159_ (.A1(_03067_),
    .A2(_04013_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09160_ (.I(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09161_ (.I(_04103_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09162_ (.A1(\u_cpu.rf_ram.memory[128][0] ),
    .A2(_04105_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09163_ (.A1(_04083_),
    .A2(_04104_),
    .B(_04106_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09164_ (.A1(\u_cpu.rf_ram.memory[128][1] ),
    .A2(_04105_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09165_ (.A1(_04088_),
    .A2(_04104_),
    .B(_04107_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09166_ (.I(_04103_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09167_ (.A1(\u_cpu.rf_ram.memory[128][2] ),
    .A2(_04108_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09168_ (.A1(_04090_),
    .A2(_04104_),
    .B(_04109_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09169_ (.A1(\u_cpu.rf_ram.memory[128][3] ),
    .A2(_04108_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09170_ (.A1(_04093_),
    .A2(_04104_),
    .B(_04110_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09171_ (.A1(\u_cpu.rf_ram.memory[128][4] ),
    .A2(_04108_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09172_ (.A1(_04095_),
    .A2(_04104_),
    .B(_04111_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09173_ (.A1(\u_cpu.rf_ram.memory[128][5] ),
    .A2(_04108_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09174_ (.A1(_04097_),
    .A2(_04105_),
    .B(_04112_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09175_ (.A1(\u_cpu.rf_ram.memory[128][6] ),
    .A2(_04108_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09176_ (.A1(_04099_),
    .A2(_04105_),
    .B(_04113_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09177_ (.A1(\u_cpu.rf_ram.memory[128][7] ),
    .A2(_04103_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09178_ (.A1(_04101_),
    .A2(_04105_),
    .B(_04114_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09179_ (.A1(_03230_),
    .A2(_03356_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09180_ (.I(_04115_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09181_ (.I(_04115_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09182_ (.A1(\u_cpu.rf_ram.memory[127][0] ),
    .A2(_04117_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09183_ (.A1(_04083_),
    .A2(_04116_),
    .B(_04118_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09184_ (.A1(\u_cpu.rf_ram.memory[127][1] ),
    .A2(_04117_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09185_ (.A1(_04088_),
    .A2(_04116_),
    .B(_04119_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09186_ (.I(_04115_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09187_ (.A1(\u_cpu.rf_ram.memory[127][2] ),
    .A2(_04120_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09188_ (.A1(_04090_),
    .A2(_04116_),
    .B(_04121_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09189_ (.A1(\u_cpu.rf_ram.memory[127][3] ),
    .A2(_04120_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09190_ (.A1(_04093_),
    .A2(_04116_),
    .B(_04122_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09191_ (.A1(\u_cpu.rf_ram.memory[127][4] ),
    .A2(_04120_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09192_ (.A1(_04095_),
    .A2(_04116_),
    .B(_04123_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(\u_cpu.rf_ram.memory[127][5] ),
    .A2(_04120_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09194_ (.A1(_04097_),
    .A2(_04117_),
    .B(_04124_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(\u_cpu.rf_ram.memory[127][6] ),
    .A2(_04120_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09196_ (.A1(_04099_),
    .A2(_04117_),
    .B(_04125_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09197_ (.A1(\u_cpu.rf_ram.memory[127][7] ),
    .A2(_04115_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09198_ (.A1(_04101_),
    .A2(_04117_),
    .B(_04126_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09199_ (.A1(_03082_),
    .A2(_03356_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09200_ (.I(_04127_),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09201_ (.I(_04127_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09202_ (.A1(\u_cpu.rf_ram.memory[126][0] ),
    .A2(_04129_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09203_ (.A1(_04083_),
    .A2(_04128_),
    .B(_04130_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09204_ (.A1(\u_cpu.rf_ram.memory[126][1] ),
    .A2(_04129_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09205_ (.A1(_04088_),
    .A2(_04128_),
    .B(_04131_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09206_ (.I(_04127_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09207_ (.A1(\u_cpu.rf_ram.memory[126][2] ),
    .A2(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09208_ (.A1(_04090_),
    .A2(_04128_),
    .B(_04133_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09209_ (.A1(\u_cpu.rf_ram.memory[126][3] ),
    .A2(_04132_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09210_ (.A1(_04093_),
    .A2(_04128_),
    .B(_04134_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09211_ (.A1(\u_cpu.rf_ram.memory[126][4] ),
    .A2(_04132_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09212_ (.A1(_04095_),
    .A2(_04128_),
    .B(_04135_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09213_ (.A1(\u_cpu.rf_ram.memory[126][5] ),
    .A2(_04132_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09214_ (.A1(_04097_),
    .A2(_04129_),
    .B(_04136_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(\u_cpu.rf_ram.memory[126][6] ),
    .A2(_04132_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09216_ (.A1(_04099_),
    .A2(_04129_),
    .B(_04137_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09217_ (.A1(\u_cpu.rf_ram.memory[126][7] ),
    .A2(_04127_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09218_ (.A1(_04101_),
    .A2(_04129_),
    .B(_04138_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09219_ (.A1(_03131_),
    .A2(_03356_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09220_ (.I(_04139_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09221_ (.I(_04139_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09222_ (.A1(\u_cpu.rf_ram.memory[125][0] ),
    .A2(_04141_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09223_ (.A1(_04083_),
    .A2(_04140_),
    .B(_04142_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09224_ (.A1(\u_cpu.rf_ram.memory[125][1] ),
    .A2(_04141_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09225_ (.A1(_04088_),
    .A2(_04140_),
    .B(_04143_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09226_ (.I(_04139_),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09227_ (.A1(\u_cpu.rf_ram.memory[125][2] ),
    .A2(_04144_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09228_ (.A1(_04090_),
    .A2(_04140_),
    .B(_04145_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09229_ (.A1(\u_cpu.rf_ram.memory[125][3] ),
    .A2(_04144_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09230_ (.A1(_04093_),
    .A2(_04140_),
    .B(_04146_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09231_ (.A1(\u_cpu.rf_ram.memory[125][4] ),
    .A2(_04144_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09232_ (.A1(_04095_),
    .A2(_04140_),
    .B(_04147_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(\u_cpu.rf_ram.memory[125][5] ),
    .A2(_04144_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09234_ (.A1(_04097_),
    .A2(_04141_),
    .B(_04148_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09235_ (.A1(\u_cpu.rf_ram.memory[125][6] ),
    .A2(_04144_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09236_ (.A1(_04099_),
    .A2(_04141_),
    .B(_04149_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09237_ (.A1(\u_cpu.rf_ram.memory[125][7] ),
    .A2(_04139_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09238_ (.A1(_04101_),
    .A2(_04141_),
    .B(_04150_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09239_ (.I(_02905_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09240_ (.I(_04151_),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09241_ (.A1(_03152_),
    .A2(_03356_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09242_ (.I(_04153_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09243_ (.I(_04153_),
    .Z(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09244_ (.A1(\u_cpu.rf_ram.memory[124][0] ),
    .A2(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09245_ (.A1(_04152_),
    .A2(_04154_),
    .B(_04156_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09246_ (.I(_02912_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09247_ (.I(_04157_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09248_ (.A1(\u_cpu.rf_ram.memory[124][1] ),
    .A2(_04155_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09249_ (.A1(_04158_),
    .A2(_04154_),
    .B(_04159_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09250_ (.I(_02918_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09251_ (.I(_04160_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09252_ (.I(_04153_),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09253_ (.A1(\u_cpu.rf_ram.memory[124][2] ),
    .A2(_04162_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09254_ (.A1(_04161_),
    .A2(_04154_),
    .B(_04163_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09255_ (.I(_02925_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09256_ (.I(_04164_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09257_ (.A1(\u_cpu.rf_ram.memory[124][3] ),
    .A2(_04162_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09258_ (.A1(_04165_),
    .A2(_04154_),
    .B(_04166_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09259_ (.I(_02931_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09260_ (.I(_04167_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09261_ (.A1(\u_cpu.rf_ram.memory[124][4] ),
    .A2(_04162_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09262_ (.A1(_04168_),
    .A2(_04154_),
    .B(_04169_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09263_ (.I(_02937_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09264_ (.I(_04170_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09265_ (.A1(\u_cpu.rf_ram.memory[124][5] ),
    .A2(_04162_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09266_ (.A1(_04171_),
    .A2(_04155_),
    .B(_04172_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09267_ (.I(_02943_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09268_ (.I(_04173_),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09269_ (.A1(\u_cpu.rf_ram.memory[124][6] ),
    .A2(_04162_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09270_ (.A1(_04174_),
    .A2(_04155_),
    .B(_04175_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09271_ (.I(_02949_),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09272_ (.I(_04176_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09273_ (.A1(\u_cpu.rf_ram.memory[124][7] ),
    .A2(_04153_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09274_ (.A1(_04177_),
    .A2(_04155_),
    .B(_04178_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09275_ (.I(_03355_),
    .Z(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09276_ (.A1(_03196_),
    .A2(_04179_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09277_ (.I(_04180_),
    .Z(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09278_ (.I(_04180_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09279_ (.A1(\u_cpu.rf_ram.memory[123][0] ),
    .A2(_04182_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09280_ (.A1(_04152_),
    .A2(_04181_),
    .B(_04183_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09281_ (.A1(\u_cpu.rf_ram.memory[123][1] ),
    .A2(_04182_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09282_ (.A1(_04158_),
    .A2(_04181_),
    .B(_04184_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09283_ (.I(_04180_),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09284_ (.A1(\u_cpu.rf_ram.memory[123][2] ),
    .A2(_04185_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09285_ (.A1(_04161_),
    .A2(_04181_),
    .B(_04186_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09286_ (.A1(\u_cpu.rf_ram.memory[123][3] ),
    .A2(_04185_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09287_ (.A1(_04165_),
    .A2(_04181_),
    .B(_04187_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09288_ (.A1(\u_cpu.rf_ram.memory[123][4] ),
    .A2(_04185_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09289_ (.A1(_04168_),
    .A2(_04181_),
    .B(_04188_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09290_ (.A1(\u_cpu.rf_ram.memory[123][5] ),
    .A2(_04185_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09291_ (.A1(_04171_),
    .A2(_04182_),
    .B(_04189_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09292_ (.A1(\u_cpu.rf_ram.memory[123][6] ),
    .A2(_04185_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09293_ (.A1(_04174_),
    .A2(_04182_),
    .B(_04190_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09294_ (.A1(\u_cpu.rf_ram.memory[123][7] ),
    .A2(_04180_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09295_ (.A1(_04177_),
    .A2(_04182_),
    .B(_04191_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(_03181_),
    .A2(_03453_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09297_ (.I(_04192_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09298_ (.I(_04192_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09299_ (.A1(\u_cpu.rf_ram.memory[38][0] ),
    .A2(_04194_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09300_ (.A1(_04152_),
    .A2(_04193_),
    .B(_04195_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09301_ (.A1(\u_cpu.rf_ram.memory[38][1] ),
    .A2(_04194_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09302_ (.A1(_04158_),
    .A2(_04193_),
    .B(_04196_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09303_ (.I(_04192_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09304_ (.A1(\u_cpu.rf_ram.memory[38][2] ),
    .A2(_04197_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09305_ (.A1(_04161_),
    .A2(_04193_),
    .B(_04198_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09306_ (.A1(\u_cpu.rf_ram.memory[38][3] ),
    .A2(_04197_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09307_ (.A1(_04165_),
    .A2(_04193_),
    .B(_04199_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09308_ (.A1(\u_cpu.rf_ram.memory[38][4] ),
    .A2(_04197_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09309_ (.A1(_04168_),
    .A2(_04193_),
    .B(_04200_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09310_ (.A1(\u_cpu.rf_ram.memory[38][5] ),
    .A2(_04197_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09311_ (.A1(_04171_),
    .A2(_04194_),
    .B(_04201_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09312_ (.A1(\u_cpu.rf_ram.memory[38][6] ),
    .A2(_04197_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09313_ (.A1(_04174_),
    .A2(_04194_),
    .B(_04202_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09314_ (.A1(\u_cpu.rf_ram.memory[38][7] ),
    .A2(_04192_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09315_ (.A1(_04177_),
    .A2(_04194_),
    .B(_04203_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09316_ (.A1(_02960_),
    .A2(_03104_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09317_ (.I(_04204_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09318_ (.I(_04204_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09319_ (.A1(\u_cpu.rf_ram.memory[37][0] ),
    .A2(_04206_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09320_ (.A1(_04152_),
    .A2(_04205_),
    .B(_04207_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09321_ (.A1(\u_cpu.rf_ram.memory[37][1] ),
    .A2(_04206_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09322_ (.A1(_04158_),
    .A2(_04205_),
    .B(_04208_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09323_ (.I(_04204_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09324_ (.A1(\u_cpu.rf_ram.memory[37][2] ),
    .A2(_04209_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09325_ (.A1(_04161_),
    .A2(_04205_),
    .B(_04210_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09326_ (.A1(\u_cpu.rf_ram.memory[37][3] ),
    .A2(_04209_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09327_ (.A1(_04165_),
    .A2(_04205_),
    .B(_04211_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(\u_cpu.rf_ram.memory[37][4] ),
    .A2(_04209_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09329_ (.A1(_04168_),
    .A2(_04205_),
    .B(_04212_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09330_ (.A1(\u_cpu.rf_ram.memory[37][5] ),
    .A2(_04209_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09331_ (.A1(_04171_),
    .A2(_04206_),
    .B(_04213_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09332_ (.A1(\u_cpu.rf_ram.memory[37][6] ),
    .A2(_04209_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09333_ (.A1(_04174_),
    .A2(_04206_),
    .B(_04214_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09334_ (.A1(\u_cpu.rf_ram.memory[37][7] ),
    .A2(_04204_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09335_ (.A1(_04177_),
    .A2(_04206_),
    .B(_04215_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09336_ (.A1(_03012_),
    .A2(_03104_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09337_ (.I(_04216_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09338_ (.I(_04216_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09339_ (.A1(\u_cpu.rf_ram.memory[36][0] ),
    .A2(_04218_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09340_ (.A1(_04152_),
    .A2(_04217_),
    .B(_04219_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09341_ (.A1(\u_cpu.rf_ram.memory[36][1] ),
    .A2(_04218_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09342_ (.A1(_04158_),
    .A2(_04217_),
    .B(_04220_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09343_ (.I(_04216_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09344_ (.A1(\u_cpu.rf_ram.memory[36][2] ),
    .A2(_04221_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09345_ (.A1(_04161_),
    .A2(_04217_),
    .B(_04222_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09346_ (.A1(\u_cpu.rf_ram.memory[36][3] ),
    .A2(_04221_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09347_ (.A1(_04165_),
    .A2(_04217_),
    .B(_04223_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09348_ (.A1(\u_cpu.rf_ram.memory[36][4] ),
    .A2(_04221_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09349_ (.A1(_04168_),
    .A2(_04217_),
    .B(_04224_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09350_ (.A1(\u_cpu.rf_ram.memory[36][5] ),
    .A2(_04221_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09351_ (.A1(_04171_),
    .A2(_04218_),
    .B(_04225_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09352_ (.A1(\u_cpu.rf_ram.memory[36][6] ),
    .A2(_04221_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09353_ (.A1(_04174_),
    .A2(_04218_),
    .B(_04226_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09354_ (.A1(\u_cpu.rf_ram.memory[36][7] ),
    .A2(_04216_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09355_ (.A1(_04177_),
    .A2(_04218_),
    .B(_04227_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09356_ (.I(_02505_),
    .Z(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09357_ (.A1(_04228_),
    .A2(_03281_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09358_ (.A1(_03270_),
    .A2(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09359_ (.I(_04230_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09360_ (.A1(_02498_),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09361_ (.A1(_02498_),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09362_ (.A1(_03271_),
    .A2(_04231_),
    .A3(_04232_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09363_ (.I(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09364_ (.I(_02621_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09365_ (.A1(_04233_),
    .A2(_04232_),
    .B(_04234_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09366_ (.A1(_04233_),
    .A2(_04232_),
    .B(_04235_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09367_ (.I(\u_cpu.cpu.mem_bytecnt[1] ),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09368_ (.A1(_04233_),
    .A2(_04232_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09369_ (.A1(_04236_),
    .A2(_04237_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09370_ (.A1(_03272_),
    .A2(_04238_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09371_ (.I(\u_cpu.rf_ram_if.rgnt ),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09372_ (.A1(_04239_),
    .A2(_03294_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09373_ (.A1(_03270_),
    .A2(_04228_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09374_ (.I(_04241_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09375_ (.A1(_02498_),
    .A2(_04242_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09376_ (.A1(_03271_),
    .A2(_02462_),
    .A3(_04240_),
    .B(_04243_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09377_ (.A1(_04234_),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09378_ (.I(_04244_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09379_ (.A1(_03272_),
    .A2(_02573_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09380_ (.A1(_04234_),
    .A2(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09381_ (.I(_04245_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09382_ (.I(_04151_),
    .Z(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09383_ (.A1(_02899_),
    .A2(_03197_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09384_ (.I(_04247_),
    .Z(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09385_ (.I(_04247_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09386_ (.A1(\u_cpu.rf_ram.memory[91][0] ),
    .A2(_04249_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09387_ (.A1(_04246_),
    .A2(_04248_),
    .B(_04250_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09388_ (.I(_04157_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09389_ (.A1(\u_cpu.rf_ram.memory[91][1] ),
    .A2(_04249_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09390_ (.A1(_04251_),
    .A2(_04248_),
    .B(_04252_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09391_ (.I(_04160_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09392_ (.I(_04247_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09393_ (.A1(\u_cpu.rf_ram.memory[91][2] ),
    .A2(_04254_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09394_ (.A1(_04253_),
    .A2(_04248_),
    .B(_04255_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09395_ (.I(_04164_),
    .Z(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09396_ (.A1(\u_cpu.rf_ram.memory[91][3] ),
    .A2(_04254_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09397_ (.A1(_04256_),
    .A2(_04248_),
    .B(_04257_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09398_ (.I(_04167_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09399_ (.A1(\u_cpu.rf_ram.memory[91][4] ),
    .A2(_04254_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09400_ (.A1(_04258_),
    .A2(_04248_),
    .B(_04259_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09401_ (.I(_04170_),
    .Z(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09402_ (.A1(\u_cpu.rf_ram.memory[91][5] ),
    .A2(_04254_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09403_ (.A1(_04260_),
    .A2(_04249_),
    .B(_04261_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09404_ (.I(_04173_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09405_ (.A1(\u_cpu.rf_ram.memory[91][6] ),
    .A2(_04254_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09406_ (.A1(_04262_),
    .A2(_04249_),
    .B(_04263_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09407_ (.I(_04176_),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09408_ (.A1(\u_cpu.rf_ram.memory[91][7] ),
    .A2(_04247_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09409_ (.A1(_04264_),
    .A2(_04249_),
    .B(_04265_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09410_ (.A1(_02899_),
    .A2(_03102_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09411_ (.I(_04266_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09412_ (.I(_04266_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09413_ (.A1(\u_cpu.rf_ram.memory[90][0] ),
    .A2(_04268_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09414_ (.A1(_04246_),
    .A2(_04267_),
    .B(_04269_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09415_ (.A1(\u_cpu.rf_ram.memory[90][1] ),
    .A2(_04268_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09416_ (.A1(_04251_),
    .A2(_04267_),
    .B(_04270_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09417_ (.I(_04266_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09418_ (.A1(\u_cpu.rf_ram.memory[90][2] ),
    .A2(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09419_ (.A1(_04253_),
    .A2(_04267_),
    .B(_04272_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09420_ (.A1(\u_cpu.rf_ram.memory[90][3] ),
    .A2(_04271_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09421_ (.A1(_04256_),
    .A2(_04267_),
    .B(_04273_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09422_ (.A1(\u_cpu.rf_ram.memory[90][4] ),
    .A2(_04271_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09423_ (.A1(_04258_),
    .A2(_04267_),
    .B(_04274_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09424_ (.A1(\u_cpu.rf_ram.memory[90][5] ),
    .A2(_04271_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09425_ (.A1(_04260_),
    .A2(_04268_),
    .B(_04275_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09426_ (.A1(\u_cpu.rf_ram.memory[90][6] ),
    .A2(_04271_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09427_ (.A1(_04262_),
    .A2(_04268_),
    .B(_04276_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09428_ (.A1(\u_cpu.rf_ram.memory[90][7] ),
    .A2(_04266_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09429_ (.A1(_04264_),
    .A2(_04268_),
    .B(_04277_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09430_ (.A1(_02614_),
    .A2(_02616_),
    .A3(_02613_),
    .Z(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09431_ (.A1(_03273_),
    .A2(_04242_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09432_ (.A1(_03271_),
    .A2(_04229_),
    .A3(_04278_),
    .B(_04279_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09433_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_04242_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09434_ (.I(_02558_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09435_ (.A1(_02492_),
    .A2(_02487_),
    .B(_02485_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09436_ (.A1(_02480_),
    .A2(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09437_ (.A1(_02478_),
    .A2(_04282_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09438_ (.A1(_02482_),
    .A2(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09439_ (.A1(_04283_),
    .A2(_04285_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09440_ (.A1(_02491_),
    .A2(_02522_),
    .B1(_04283_),
    .B2(_04285_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09441_ (.I(\u_cpu.cpu.alu.cmp_r ),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09442_ (.A1(_04288_),
    .A2(_02548_),
    .B(_02495_),
    .C(_02487_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09443_ (.A1(_04286_),
    .A2(_04287_),
    .B1(_04289_),
    .B2(_02563_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09444_ (.A1(_02493_),
    .A2(_04290_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09445_ (.A1(_04281_),
    .A2(_04291_),
    .B(_00773_),
    .C(_02617_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09446_ (.A1(_04280_),
    .A2(_04292_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09447_ (.A1(_04236_),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(_04233_),
    .A4(_00780_),
    .Z(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09448_ (.I(_04293_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09449_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_04242_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09450_ (.A1(_03272_),
    .A2(_04229_),
    .B(_04294_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09451_ (.I(_02898_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09452_ (.A1(_04295_),
    .A2(_03153_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09453_ (.I(_04296_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09454_ (.I(_04296_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09455_ (.A1(\u_cpu.rf_ram.memory[92][0] ),
    .A2(_04298_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09456_ (.A1(_04246_),
    .A2(_04297_),
    .B(_04299_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09457_ (.A1(\u_cpu.rf_ram.memory[92][1] ),
    .A2(_04298_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09458_ (.A1(_04251_),
    .A2(_04297_),
    .B(_04300_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09459_ (.I(_04296_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(\u_cpu.rf_ram.memory[92][2] ),
    .A2(_04301_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09461_ (.A1(_04253_),
    .A2(_04297_),
    .B(_04302_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09462_ (.A1(\u_cpu.rf_ram.memory[92][3] ),
    .A2(_04301_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09463_ (.A1(_04256_),
    .A2(_04297_),
    .B(_04303_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09464_ (.A1(\u_cpu.rf_ram.memory[92][4] ),
    .A2(_04301_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09465_ (.A1(_04258_),
    .A2(_04297_),
    .B(_04304_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09466_ (.A1(\u_cpu.rf_ram.memory[92][5] ),
    .A2(_04301_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09467_ (.A1(_04260_),
    .A2(_04298_),
    .B(_04305_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09468_ (.A1(\u_cpu.rf_ram.memory[92][6] ),
    .A2(_04301_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09469_ (.A1(_04262_),
    .A2(_04298_),
    .B(_04306_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09470_ (.A1(\u_cpu.rf_ram.memory[92][7] ),
    .A2(_04296_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09471_ (.A1(_04264_),
    .A2(_04298_),
    .B(_04307_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09472_ (.A1(_03103_),
    .A2(_03480_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09473_ (.I(_04308_),
    .Z(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09474_ (.I(_04308_),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09475_ (.A1(\u_cpu.rf_ram.memory[35][0] ),
    .A2(_04310_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09476_ (.A1(_04246_),
    .A2(_04309_),
    .B(_04311_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09477_ (.A1(\u_cpu.rf_ram.memory[35][1] ),
    .A2(_04310_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09478_ (.A1(_04251_),
    .A2(_04309_),
    .B(_04312_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09479_ (.I(_04308_),
    .Z(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09480_ (.A1(\u_cpu.rf_ram.memory[35][2] ),
    .A2(_04313_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09481_ (.A1(_04253_),
    .A2(_04309_),
    .B(_04314_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09482_ (.A1(\u_cpu.rf_ram.memory[35][3] ),
    .A2(_04313_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09483_ (.A1(_04256_),
    .A2(_04309_),
    .B(_04315_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(\u_cpu.rf_ram.memory[35][4] ),
    .A2(_04313_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09485_ (.A1(_04258_),
    .A2(_04309_),
    .B(_04316_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09486_ (.A1(\u_cpu.rf_ram.memory[35][5] ),
    .A2(_04313_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09487_ (.A1(_04260_),
    .A2(_04310_),
    .B(_04317_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09488_ (.A1(\u_cpu.rf_ram.memory[35][6] ),
    .A2(_04313_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09489_ (.A1(_04262_),
    .A2(_04310_),
    .B(_04318_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(\u_cpu.rf_ram.memory[35][7] ),
    .A2(_04308_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09491_ (.A1(_04264_),
    .A2(_04310_),
    .B(_04319_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09492_ (.A1(_02890_),
    .A2(_03130_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09493_ (.I(_04320_),
    .Z(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09494_ (.I(_04320_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09495_ (.A1(\u_cpu.rf_ram.memory[34][0] ),
    .A2(_04322_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09496_ (.A1(_04246_),
    .A2(_04321_),
    .B(_04323_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09497_ (.A1(\u_cpu.rf_ram.memory[34][1] ),
    .A2(_04322_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09498_ (.A1(_04251_),
    .A2(_04321_),
    .B(_04324_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09499_ (.I(_04320_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09500_ (.A1(\u_cpu.rf_ram.memory[34][2] ),
    .A2(_04325_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09501_ (.A1(_04253_),
    .A2(_04321_),
    .B(_04326_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09502_ (.A1(\u_cpu.rf_ram.memory[34][3] ),
    .A2(_04325_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09503_ (.A1(_04256_),
    .A2(_04321_),
    .B(_04327_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09504_ (.A1(\u_cpu.rf_ram.memory[34][4] ),
    .A2(_04325_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09505_ (.A1(_04258_),
    .A2(_04321_),
    .B(_04328_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09506_ (.A1(\u_cpu.rf_ram.memory[34][5] ),
    .A2(_04325_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09507_ (.A1(_04260_),
    .A2(_04322_),
    .B(_04329_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09508_ (.A1(\u_cpu.rf_ram.memory[34][6] ),
    .A2(_04325_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09509_ (.A1(_04262_),
    .A2(_04322_),
    .B(_04330_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09510_ (.A1(\u_cpu.rf_ram.memory[34][7] ),
    .A2(_04320_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09511_ (.A1(_04264_),
    .A2(_04322_),
    .B(_04331_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09512_ (.I(_04151_),
    .Z(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09513_ (.A1(_02960_),
    .A2(_04179_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09514_ (.I(_04333_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09515_ (.I(_04333_),
    .Z(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09516_ (.A1(\u_cpu.rf_ram.memory[117][0] ),
    .A2(_04335_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09517_ (.A1(_04332_),
    .A2(_04334_),
    .B(_04336_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09518_ (.I(_04157_),
    .Z(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09519_ (.A1(\u_cpu.rf_ram.memory[117][1] ),
    .A2(_04335_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09520_ (.A1(_04337_),
    .A2(_04334_),
    .B(_04338_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09521_ (.I(_04160_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09522_ (.I(_04333_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09523_ (.A1(\u_cpu.rf_ram.memory[117][2] ),
    .A2(_04340_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09524_ (.A1(_04339_),
    .A2(_04334_),
    .B(_04341_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09525_ (.I(_04164_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09526_ (.A1(\u_cpu.rf_ram.memory[117][3] ),
    .A2(_04340_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09527_ (.A1(_04342_),
    .A2(_04334_),
    .B(_04343_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09528_ (.I(_04167_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09529_ (.A1(\u_cpu.rf_ram.memory[117][4] ),
    .A2(_04340_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09530_ (.A1(_04344_),
    .A2(_04334_),
    .B(_04345_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09531_ (.I(_04170_),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09532_ (.A1(\u_cpu.rf_ram.memory[117][5] ),
    .A2(_04340_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09533_ (.A1(_04346_),
    .A2(_04335_),
    .B(_04347_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09534_ (.I(_04173_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09535_ (.A1(\u_cpu.rf_ram.memory[117][6] ),
    .A2(_04340_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09536_ (.A1(_04348_),
    .A2(_04335_),
    .B(_04349_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09537_ (.I(_04176_),
    .Z(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09538_ (.A1(\u_cpu.rf_ram.memory[117][7] ),
    .A2(_04333_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09539_ (.A1(_04350_),
    .A2(_04335_),
    .B(_04351_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09540_ (.A1(_03327_),
    .A2(_04179_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09541_ (.I(_04352_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09542_ (.I(_04352_),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09543_ (.A1(\u_cpu.rf_ram.memory[120][0] ),
    .A2(_04354_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09544_ (.A1(_04332_),
    .A2(_04353_),
    .B(_04355_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09545_ (.A1(\u_cpu.rf_ram.memory[120][1] ),
    .A2(_04354_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09546_ (.A1(_04337_),
    .A2(_04353_),
    .B(_04356_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09547_ (.I(_04352_),
    .Z(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09548_ (.A1(\u_cpu.rf_ram.memory[120][2] ),
    .A2(_04357_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09549_ (.A1(_04339_),
    .A2(_04353_),
    .B(_04358_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09550_ (.A1(\u_cpu.rf_ram.memory[120][3] ),
    .A2(_04357_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09551_ (.A1(_04342_),
    .A2(_04353_),
    .B(_04359_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09552_ (.A1(\u_cpu.rf_ram.memory[120][4] ),
    .A2(_04357_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09553_ (.A1(_04344_),
    .A2(_04353_),
    .B(_04360_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09554_ (.A1(\u_cpu.rf_ram.memory[120][5] ),
    .A2(_04357_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09555_ (.A1(_04346_),
    .A2(_04354_),
    .B(_04361_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09556_ (.A1(\u_cpu.rf_ram.memory[120][6] ),
    .A2(_04357_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09557_ (.A1(_04348_),
    .A2(_04354_),
    .B(_04362_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09558_ (.A1(\u_cpu.rf_ram.memory[120][7] ),
    .A2(_04352_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09559_ (.A1(_04350_),
    .A2(_04354_),
    .B(_04363_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09560_ (.A1(_03355_),
    .A2(_03453_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09561_ (.I(_04364_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09562_ (.I(_04364_),
    .Z(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09563_ (.A1(\u_cpu.rf_ram.memory[118][0] ),
    .A2(_04366_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09564_ (.A1(_04332_),
    .A2(_04365_),
    .B(_04367_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09565_ (.A1(\u_cpu.rf_ram.memory[118][1] ),
    .A2(_04366_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09566_ (.A1(_04337_),
    .A2(_04365_),
    .B(_04368_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09567_ (.I(_04364_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09568_ (.A1(\u_cpu.rf_ram.memory[118][2] ),
    .A2(_04369_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09569_ (.A1(_04339_),
    .A2(_04365_),
    .B(_04370_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09570_ (.A1(\u_cpu.rf_ram.memory[118][3] ),
    .A2(_04369_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09571_ (.A1(_04342_),
    .A2(_04365_),
    .B(_04371_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(\u_cpu.rf_ram.memory[118][4] ),
    .A2(_04369_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09573_ (.A1(_04344_),
    .A2(_04365_),
    .B(_04372_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09574_ (.A1(\u_cpu.rf_ram.memory[118][5] ),
    .A2(_04369_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09575_ (.A1(_04346_),
    .A2(_04366_),
    .B(_04373_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09576_ (.A1(\u_cpu.rf_ram.memory[118][6] ),
    .A2(_04369_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09577_ (.A1(_04348_),
    .A2(_04366_),
    .B(_04374_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09578_ (.A1(\u_cpu.rf_ram.memory[118][7] ),
    .A2(_04364_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09579_ (.A1(_04350_),
    .A2(_04366_),
    .B(_04375_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09580_ (.A1(_03182_),
    .A2(_04179_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09581_ (.I(_04376_),
    .Z(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09582_ (.I(_04376_),
    .Z(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09583_ (.A1(\u_cpu.rf_ram.memory[121][0] ),
    .A2(_04378_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09584_ (.A1(_04332_),
    .A2(_04377_),
    .B(_04379_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09585_ (.A1(\u_cpu.rf_ram.memory[121][1] ),
    .A2(_04378_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09586_ (.A1(_04337_),
    .A2(_04377_),
    .B(_04380_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09587_ (.I(_04376_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09588_ (.A1(\u_cpu.rf_ram.memory[121][2] ),
    .A2(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09589_ (.A1(_04339_),
    .A2(_04377_),
    .B(_04382_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09590_ (.A1(\u_cpu.rf_ram.memory[121][3] ),
    .A2(_04381_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09591_ (.A1(_04342_),
    .A2(_04377_),
    .B(_04383_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09592_ (.A1(\u_cpu.rf_ram.memory[121][4] ),
    .A2(_04381_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09593_ (.A1(_04344_),
    .A2(_04377_),
    .B(_04384_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09594_ (.A1(\u_cpu.rf_ram.memory[121][5] ),
    .A2(_04381_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09595_ (.A1(_04346_),
    .A2(_04378_),
    .B(_04385_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09596_ (.A1(\u_cpu.rf_ram.memory[121][6] ),
    .A2(_04381_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09597_ (.A1(_04348_),
    .A2(_04378_),
    .B(_04386_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09598_ (.A1(\u_cpu.rf_ram.memory[121][7] ),
    .A2(_04376_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09599_ (.A1(_04350_),
    .A2(_04378_),
    .B(_04387_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09600_ (.A1(_03037_),
    .A2(_03328_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09601_ (.I(_04388_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09602_ (.I(_04388_),
    .Z(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09603_ (.A1(\u_cpu.rf_ram.memory[8][0] ),
    .A2(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09604_ (.A1(_04062_),
    .A2(_04389_),
    .B(_04391_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09605_ (.A1(\u_cpu.rf_ram.memory[8][1] ),
    .A2(_04390_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09606_ (.A1(_04068_),
    .A2(_04389_),
    .B(_04392_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09607_ (.I(_04388_),
    .Z(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09608_ (.A1(\u_cpu.rf_ram.memory[8][2] ),
    .A2(_04393_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09609_ (.A1(_04070_),
    .A2(_04389_),
    .B(_04394_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09610_ (.A1(\u_cpu.rf_ram.memory[8][3] ),
    .A2(_04393_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09611_ (.A1(_04073_),
    .A2(_04389_),
    .B(_04395_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09612_ (.A1(\u_cpu.rf_ram.memory[8][4] ),
    .A2(_04393_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09613_ (.A1(_04075_),
    .A2(_04389_),
    .B(_04396_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09614_ (.A1(\u_cpu.rf_ram.memory[8][5] ),
    .A2(_04393_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09615_ (.A1(_04077_),
    .A2(_04390_),
    .B(_04397_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09616_ (.A1(\u_cpu.rf_ram.memory[8][6] ),
    .A2(_04393_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09617_ (.A1(_04079_),
    .A2(_04390_),
    .B(_04398_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09618_ (.A1(\u_cpu.rf_ram.memory[8][7] ),
    .A2(_04388_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09619_ (.A1(_04081_),
    .A2(_04390_),
    .B(_04399_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09620_ (.A1(_03256_),
    .A2(_03197_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09621_ (.I(_04400_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09622_ (.I(_04401_),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09623_ (.I(_04401_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09624_ (.A1(\u_cpu.rf_ram.memory[11][0] ),
    .A2(_04403_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09625_ (.A1(_04062_),
    .A2(_04402_),
    .B(_04404_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09626_ (.A1(\u_cpu.rf_ram.memory[11][1] ),
    .A2(_04403_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09627_ (.A1(_04068_),
    .A2(_04402_),
    .B(_04405_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09628_ (.I(_04401_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09629_ (.A1(\u_cpu.rf_ram.memory[11][2] ),
    .A2(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09630_ (.A1(_04070_),
    .A2(_04402_),
    .B(_04407_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09631_ (.A1(\u_cpu.rf_ram.memory[11][3] ),
    .A2(_04406_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09632_ (.A1(_04073_),
    .A2(_04402_),
    .B(_04408_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09633_ (.A1(\u_cpu.rf_ram.memory[11][4] ),
    .A2(_04406_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09634_ (.A1(_04075_),
    .A2(_04402_),
    .B(_04409_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09635_ (.A1(\u_cpu.rf_ram.memory[11][5] ),
    .A2(_04406_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09636_ (.A1(_04077_),
    .A2(_04403_),
    .B(_04410_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09637_ (.A1(\u_cpu.rf_ram.memory[11][6] ),
    .A2(_04406_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09638_ (.A1(_04079_),
    .A2(_04403_),
    .B(_04411_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09639_ (.A1(\u_cpu.rf_ram.memory[11][7] ),
    .A2(_04401_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09640_ (.A1(_04081_),
    .A2(_04403_),
    .B(_04412_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09641_ (.A1(_03067_),
    .A2(_04179_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09642_ (.I(_04413_),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09643_ (.I(_04413_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09644_ (.A1(\u_cpu.rf_ram.memory[112][0] ),
    .A2(_04415_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09645_ (.A1(_04332_),
    .A2(_04414_),
    .B(_04416_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09646_ (.A1(\u_cpu.rf_ram.memory[112][1] ),
    .A2(_04415_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09647_ (.A1(_04337_),
    .A2(_04414_),
    .B(_04417_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09648_ (.I(_04413_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09649_ (.A1(\u_cpu.rf_ram.memory[112][2] ),
    .A2(_04418_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09650_ (.A1(_04339_),
    .A2(_04414_),
    .B(_04419_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09651_ (.A1(\u_cpu.rf_ram.memory[112][3] ),
    .A2(_04418_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09652_ (.A1(_04342_),
    .A2(_04414_),
    .B(_04420_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09653_ (.A1(\u_cpu.rf_ram.memory[112][4] ),
    .A2(_04418_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09654_ (.A1(_04344_),
    .A2(_04414_),
    .B(_04421_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09655_ (.A1(\u_cpu.rf_ram.memory[112][5] ),
    .A2(_04418_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09656_ (.A1(_04346_),
    .A2(_04415_),
    .B(_04422_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09657_ (.A1(\u_cpu.rf_ram.memory[112][6] ),
    .A2(_04418_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09658_ (.A1(_04348_),
    .A2(_04415_),
    .B(_04423_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09659_ (.A1(\u_cpu.rf_ram.memory[112][7] ),
    .A2(_04413_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09660_ (.A1(_04350_),
    .A2(_04415_),
    .B(_04424_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09661_ (.I(_04151_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09662_ (.I(_03355_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09663_ (.A1(_03101_),
    .A2(_04426_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09664_ (.I(_04427_),
    .Z(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09665_ (.I(_04427_),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09666_ (.A1(\u_cpu.rf_ram.memory[122][0] ),
    .A2(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09667_ (.A1(_04425_),
    .A2(_04428_),
    .B(_04430_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09668_ (.I(_04157_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09669_ (.A1(\u_cpu.rf_ram.memory[122][1] ),
    .A2(_04429_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09670_ (.A1(_04431_),
    .A2(_04428_),
    .B(_04432_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09671_ (.I(_04160_),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09672_ (.I(_04427_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09673_ (.A1(\u_cpu.rf_ram.memory[122][2] ),
    .A2(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09674_ (.A1(_04433_),
    .A2(_04428_),
    .B(_04435_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09675_ (.I(_04164_),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09676_ (.A1(\u_cpu.rf_ram.memory[122][3] ),
    .A2(_04434_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09677_ (.A1(_04436_),
    .A2(_04428_),
    .B(_04437_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09678_ (.I(_04167_),
    .Z(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09679_ (.A1(\u_cpu.rf_ram.memory[122][4] ),
    .A2(_04434_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09680_ (.A1(_04438_),
    .A2(_04428_),
    .B(_04439_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09681_ (.I(_04170_),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09682_ (.A1(\u_cpu.rf_ram.memory[122][5] ),
    .A2(_04434_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09683_ (.A1(_04440_),
    .A2(_04429_),
    .B(_04441_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09684_ (.I(_04173_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09685_ (.A1(\u_cpu.rf_ram.memory[122][6] ),
    .A2(_04434_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09686_ (.A1(_04442_),
    .A2(_04429_),
    .B(_04443_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09687_ (.I(_04176_),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09688_ (.A1(\u_cpu.rf_ram.memory[122][7] ),
    .A2(_04427_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09689_ (.A1(_04444_),
    .A2(_04429_),
    .B(_04445_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09690_ (.A1(_03166_),
    .A2(_04426_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09691_ (.I(_04446_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09692_ (.I(_04446_),
    .Z(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09693_ (.A1(\u_cpu.rf_ram.memory[115][0] ),
    .A2(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09694_ (.A1(_04425_),
    .A2(_04447_),
    .B(_04449_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09695_ (.A1(\u_cpu.rf_ram.memory[115][1] ),
    .A2(_04448_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09696_ (.A1(_04431_),
    .A2(_04447_),
    .B(_04450_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09697_ (.I(_04446_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09698_ (.A1(\u_cpu.rf_ram.memory[115][2] ),
    .A2(_04451_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09699_ (.A1(_04433_),
    .A2(_04447_),
    .B(_04452_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09700_ (.A1(\u_cpu.rf_ram.memory[115][3] ),
    .A2(_04451_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09701_ (.A1(_04436_),
    .A2(_04447_),
    .B(_04453_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09702_ (.A1(\u_cpu.rf_ram.memory[115][4] ),
    .A2(_04451_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09703_ (.A1(_04438_),
    .A2(_04447_),
    .B(_04454_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09704_ (.A1(\u_cpu.rf_ram.memory[115][5] ),
    .A2(_04451_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09705_ (.A1(_04440_),
    .A2(_04448_),
    .B(_04455_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09706_ (.A1(\u_cpu.rf_ram.memory[115][6] ),
    .A2(_04451_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09707_ (.A1(_04442_),
    .A2(_04448_),
    .B(_04456_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09708_ (.A1(\u_cpu.rf_ram.memory[115][7] ),
    .A2(_04446_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09709_ (.A1(_04444_),
    .A2(_04448_),
    .B(_04457_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09710_ (.A1(_03012_),
    .A2(_04426_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09711_ (.I(_04458_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09712_ (.I(_04458_),
    .Z(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09713_ (.A1(\u_cpu.rf_ram.memory[116][0] ),
    .A2(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09714_ (.A1(_04425_),
    .A2(_04459_),
    .B(_04461_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09715_ (.A1(\u_cpu.rf_ram.memory[116][1] ),
    .A2(_04460_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09716_ (.A1(_04431_),
    .A2(_04459_),
    .B(_04462_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09717_ (.I(_04458_),
    .Z(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09718_ (.A1(\u_cpu.rf_ram.memory[116][2] ),
    .A2(_04463_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09719_ (.A1(_04433_),
    .A2(_04459_),
    .B(_04464_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09720_ (.A1(\u_cpu.rf_ram.memory[116][3] ),
    .A2(_04463_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09721_ (.A1(_04436_),
    .A2(_04459_),
    .B(_04465_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09722_ (.A1(\u_cpu.rf_ram.memory[116][4] ),
    .A2(_04463_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09723_ (.A1(_04438_),
    .A2(_04459_),
    .B(_04466_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09724_ (.A1(\u_cpu.rf_ram.memory[116][5] ),
    .A2(_04463_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09725_ (.A1(_04440_),
    .A2(_04460_),
    .B(_04467_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09726_ (.A1(\u_cpu.rf_ram.memory[116][6] ),
    .A2(_04463_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09727_ (.A1(_04442_),
    .A2(_04460_),
    .B(_04468_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09728_ (.A1(\u_cpu.rf_ram.memory[116][7] ),
    .A2(_04458_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09729_ (.A1(_04444_),
    .A2(_04460_),
    .B(_04469_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09730_ (.A1(_02984_),
    .A2(_03130_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09731_ (.I(_04470_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09732_ (.I(_04470_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09733_ (.A1(\u_cpu.rf_ram.memory[33][0] ),
    .A2(_04472_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09734_ (.A1(_04425_),
    .A2(_04471_),
    .B(_04473_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09735_ (.A1(\u_cpu.rf_ram.memory[33][1] ),
    .A2(_04472_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09736_ (.A1(_04431_),
    .A2(_04471_),
    .B(_04474_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09737_ (.I(_04470_),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09738_ (.A1(\u_cpu.rf_ram.memory[33][2] ),
    .A2(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09739_ (.A1(_04433_),
    .A2(_04471_),
    .B(_04476_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09740_ (.A1(\u_cpu.rf_ram.memory[33][3] ),
    .A2(_04475_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09741_ (.A1(_04436_),
    .A2(_04471_),
    .B(_04477_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09742_ (.A1(\u_cpu.rf_ram.memory[33][4] ),
    .A2(_04475_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09743_ (.A1(_04438_),
    .A2(_04471_),
    .B(_04478_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09744_ (.A1(\u_cpu.rf_ram.memory[33][5] ),
    .A2(_04475_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09745_ (.A1(_04440_),
    .A2(_04472_),
    .B(_04479_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09746_ (.A1(\u_cpu.rf_ram.memory[33][6] ),
    .A2(_04475_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09747_ (.A1(_04442_),
    .A2(_04472_),
    .B(_04480_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09748_ (.A1(\u_cpu.rf_ram.memory[33][7] ),
    .A2(_04470_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09749_ (.A1(_04444_),
    .A2(_04472_),
    .B(_04481_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09750_ (.A1(_04236_),
    .A2(_02611_),
    .B(\u_cpu.cpu.bufreg.lsb[0] ),
    .C(\u_cpu.cpu.mem_bytecnt[0] ),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09751_ (.A1(_04236_),
    .A2(_02611_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09752_ (.A1(_02460_),
    .A2(_04482_),
    .A3(_04483_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09753_ (.A1(_03280_),
    .A2(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09754_ (.I(_04485_),
    .Z(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09755_ (.I(_03282_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09756_ (.A1(_02649_),
    .A2(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09757_ (.A1(_04486_),
    .A2(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09758_ (.I(_03282_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09759_ (.I(_03291_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09760_ (.I(_04491_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09761_ (.A1(_02651_),
    .A2(_04490_),
    .B(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09762_ (.A1(_02632_),
    .A2(_02622_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09763_ (.I(_04494_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09764_ (.A1(_04494_),
    .A2(_04485_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09765_ (.I(_04496_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09766_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_04495_),
    .B1(_04497_),
    .B2(_02649_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09767_ (.A1(_04489_),
    .A2(_04493_),
    .B(_04498_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09768_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_04490_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09769_ (.A1(_02649_),
    .A2(_02651_),
    .B(_04487_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09770_ (.A1(_04486_),
    .A2(_04500_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09771_ (.A1(_02651_),
    .A2(_04489_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09772_ (.A1(_04499_),
    .A2(_04501_),
    .B(_04491_),
    .C(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09773_ (.A1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_04492_),
    .B(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09774_ (.I(_04504_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09775_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_04487_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09776_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_02649_),
    .A3(_02651_),
    .B(_04487_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09777_ (.A1(_04486_),
    .A2(_04506_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09778_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_04501_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09779_ (.A1(_04505_),
    .A2(_04507_),
    .B(_04491_),
    .C(_04508_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09780_ (.A1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_04492_),
    .B(_04509_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09781_ (.I(_04510_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09782_ (.I(_04494_),
    .Z(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09783_ (.I(_04511_),
    .Z(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09784_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_04487_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09785_ (.A1(_04490_),
    .A2(_03283_),
    .B(_04513_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09786_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_04507_),
    .B1(_04514_),
    .B2(_04486_),
    .C(_04511_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09787_ (.A1(_02648_),
    .A2(_04512_),
    .B(_04515_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09788_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_03283_),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09789_ (.A1(_04490_),
    .A2(_04516_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09790_ (.A1(_03291_),
    .A2(_04485_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09791_ (.I(_04518_),
    .Z(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09792_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_04490_),
    .B(_04517_),
    .C(_04519_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09793_ (.I(_04496_),
    .Z(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09794_ (.A1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_04512_),
    .B1(_04521_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09795_ (.A1(_04520_),
    .A2(_04522_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09796_ (.A1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_04512_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09797_ (.I(_04519_),
    .Z(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09798_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_04497_),
    .B1(_04524_),
    .B2(_03289_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09799_ (.A1(_04523_),
    .A2(_04525_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09800_ (.I(_04497_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09801_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09802_ (.A1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_04512_),
    .B1(_04524_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09803_ (.A1(_04527_),
    .A2(_04528_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09804_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .A2(_04526_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09805_ (.A1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .A2(_04512_),
    .B1(_04524_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09806_ (.A1(_04529_),
    .A2(_04530_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09807_ (.I(_04496_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09808_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(_04531_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09809_ (.I(_04511_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09810_ (.I(_04518_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09811_ (.A1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_04533_),
    .B1(_04534_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09812_ (.A1(_04532_),
    .A2(_04535_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09813_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .A2(_04531_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09814_ (.A1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_04533_),
    .B1(_04534_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09815_ (.A1(_04536_),
    .A2(_04537_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09816_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .A2(_04531_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09817_ (.A1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .A2(_04533_),
    .B1(_04534_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09818_ (.A1(_04538_),
    .A2(_04539_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09819_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .A2(_04531_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09820_ (.A1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_04533_),
    .B1(_04534_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09821_ (.A1(_04540_),
    .A2(_04541_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09822_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .A2(_04531_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09823_ (.A1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_04533_),
    .B1(_04534_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09824_ (.A1(_04542_),
    .A2(_04543_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09825_ (.I(_04496_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09826_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .A2(_04544_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09827_ (.I(_04494_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09828_ (.I(_04518_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09829_ (.A1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_04546_),
    .B1(_04547_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09830_ (.A1(_04545_),
    .A2(_04548_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09831_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .A2(_04544_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09832_ (.A1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .A2(_04546_),
    .B1(_04547_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09833_ (.A1(_04549_),
    .A2(_04550_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09834_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .A2(_04544_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09835_ (.A1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .A2(_04546_),
    .B1(_04547_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09836_ (.A1(_04551_),
    .A2(_04552_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09837_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .A2(_04544_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09838_ (.A1(\u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_04546_),
    .B1(_04547_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09839_ (.A1(_04553_),
    .A2(_04554_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09840_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .A2(_04544_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09841_ (.A1(\u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_04546_),
    .B1(_04547_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09842_ (.A1(_04555_),
    .A2(_04556_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09843_ (.I(_04496_),
    .Z(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09844_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .A2(_04557_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09845_ (.I(_04494_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09846_ (.I(_04518_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09847_ (.A1(\u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_04559_),
    .B1(_04560_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09848_ (.A1(_04558_),
    .A2(_04561_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09849_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(_04557_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09850_ (.A1(\u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_04559_),
    .B1(_04560_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09851_ (.A1(_04562_),
    .A2(_04563_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09852_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .A2(_04557_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09853_ (.A1(\u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_04559_),
    .B1(_04560_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09854_ (.A1(_04564_),
    .A2(_04565_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09855_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .A2(_04557_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09856_ (.A1(\u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_04559_),
    .B1(_04560_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09857_ (.A1(_04566_),
    .A2(_04567_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09858_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .A2(_04557_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09859_ (.A1(\u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_04559_),
    .B1(_04560_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09860_ (.A1(_04568_),
    .A2(_04569_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09861_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .A2(_04521_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09862_ (.A1(\u_arbiter.i_wb_cpu_rdt[23] ),
    .A2(_04495_),
    .B1(_04519_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09863_ (.A1(_04570_),
    .A2(_04571_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09864_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .A2(_04524_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09865_ (.A1(\u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_04495_),
    .B1(_04521_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09866_ (.A1(_04572_),
    .A2(_04573_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09867_ (.A1(_04491_),
    .A2(_04486_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09868_ (.A1(\u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_04511_),
    .B1(_04497_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09869_ (.A1(_02683_),
    .A2(_04574_),
    .B(_04575_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09870_ (.A1(\u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_04492_),
    .B1(_04574_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09871_ (.A1(_02683_),
    .A2(_04526_),
    .B(_04576_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09872_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .A2(_04521_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09873_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_04495_),
    .B1(_04519_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09874_ (.A1(_04577_),
    .A2(_04578_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09875_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .A2(_04521_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09876_ (.A1(\u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_04495_),
    .B1(_04519_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09877_ (.A1(_04579_),
    .A2(_04580_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09878_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_04511_),
    .B1(_04497_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09879_ (.A1(_02690_),
    .A2(_04574_),
    .B(_04581_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09880_ (.A1(\u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_04491_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09881_ (.A1(_02690_),
    .A2(_04526_),
    .B1(_04524_),
    .B2(_02692_),
    .C(_04582_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09882_ (.A1(\u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_04492_),
    .B1(_04574_),
    .B2(_02478_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09883_ (.A1(_02692_),
    .A2(_04526_),
    .B(_04583_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09884_ (.A1(_02984_),
    .A2(_04426_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09885_ (.I(_04584_),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09886_ (.I(_04584_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09887_ (.A1(\u_cpu.rf_ram.memory[113][0] ),
    .A2(_04586_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09888_ (.A1(_04425_),
    .A2(_04585_),
    .B(_04587_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09889_ (.A1(\u_cpu.rf_ram.memory[113][1] ),
    .A2(_04586_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09890_ (.A1(_04431_),
    .A2(_04585_),
    .B(_04588_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09891_ (.I(_04584_),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09892_ (.A1(\u_cpu.rf_ram.memory[113][2] ),
    .A2(_04589_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09893_ (.A1(_04433_),
    .A2(_04585_),
    .B(_04590_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09894_ (.A1(\u_cpu.rf_ram.memory[113][3] ),
    .A2(_04589_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09895_ (.A1(_04436_),
    .A2(_04585_),
    .B(_04591_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09896_ (.A1(\u_cpu.rf_ram.memory[113][4] ),
    .A2(_04589_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09897_ (.A1(_04438_),
    .A2(_04585_),
    .B(_04592_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09898_ (.A1(\u_cpu.rf_ram.memory[113][5] ),
    .A2(_04589_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09899_ (.A1(_04440_),
    .A2(_04586_),
    .B(_04593_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09900_ (.A1(\u_cpu.rf_ram.memory[113][6] ),
    .A2(_04589_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09901_ (.A1(_04442_),
    .A2(_04586_),
    .B(_04594_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09902_ (.A1(\u_cpu.rf_ram.memory[113][7] ),
    .A2(_04584_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09903_ (.A1(_04444_),
    .A2(_04586_),
    .B(_04595_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09904_ (.I(_03275_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09905_ (.A1(_04596_),
    .A2(_02699_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09906_ (.A1(_02632_),
    .A2(_02702_),
    .A3(_04597_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09907_ (.I(_04598_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09908_ (.I(_04599_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09909_ (.I(_04600_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09910_ (.I(_02706_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09911_ (.I(_02726_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09912_ (.I(_04603_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09913_ (.I(_04604_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09914_ (.A1(_04605_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09915_ (.A1(_04602_),
    .A2(_02646_),
    .B(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09916_ (.I(_04607_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09917_ (.I0(\u_arbiter.i_wb_cpu_rdt[0] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_04604_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09918_ (.A1(_02706_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09919_ (.A1(_02706_),
    .A2(_02642_),
    .B(_04610_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09920_ (.A1(_04609_),
    .A2(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09921_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_02705_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09922_ (.A1(_04603_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09923_ (.A1(_03274_),
    .A2(\u_arbiter.i_wb_cpu_rdt[15] ),
    .B(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09924_ (.A1(_04613_),
    .A2(_04615_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09925_ (.A1(_04609_),
    .A2(_04611_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09926_ (.A1(_04616_),
    .A2(_04617_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09927_ (.A1(_04612_),
    .A2(_04618_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09928_ (.I(_04619_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09929_ (.A1(_04605_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09930_ (.A1(_03275_),
    .A2(\u_arbiter.i_wb_cpu_rdt[0] ),
    .B(_04621_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09931_ (.I(_04611_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09932_ (.A1(_04622_),
    .A2(_04623_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09933_ (.I(_04624_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09934_ (.A1(_02705_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09935_ (.A1(_03274_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_04626_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09936_ (.A1(_04613_),
    .A2(_04627_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09937_ (.I(_04628_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09938_ (.I(_04615_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09939_ (.A1(_04613_),
    .A2(_04630_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09940_ (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09941_ (.A1(_04603_),
    .A2(\u_arbiter.i_wb_cpu_rdt[11] ),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09942_ (.A1(_02705_),
    .A2(_04632_),
    .B(_04633_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09943_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_02726_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09944_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_02726_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09945_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_04603_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _09946_ (.A1(_04634_),
    .A2(_04635_),
    .A3(_04636_),
    .A4(_04637_),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09947_ (.A1(_02705_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09948_ (.A1(_03274_),
    .A2(\u_arbiter.i_wb_cpu_rdt[8] ),
    .B(_04639_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09949_ (.A1(_04638_),
    .A2(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09950_ (.A1(_04627_),
    .A2(_04631_),
    .A3(_04641_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09951_ (.A1(_04629_),
    .A2(_04642_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09952_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_04605_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09953_ (.I(_04644_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09954_ (.A1(_04638_),
    .A2(_04645_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09955_ (.A1(_04602_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09956_ (.A1(_03275_),
    .A2(\u_arbiter.i_wb_cpu_rdt[12] ),
    .B(_04647_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09957_ (.A1(_04646_),
    .A2(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09958_ (.I(_04609_),
    .Z(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09959_ (.A1(_04602_),
    .A2(_02642_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09960_ (.A1(_02707_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .B(_04651_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09961_ (.I(_04652_),
    .Z(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09962_ (.A1(_04650_),
    .A2(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09963_ (.I(_04613_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09964_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_04604_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09965_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_04604_),
    .Z(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09966_ (.A1(_04656_),
    .A2(_04657_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09967_ (.A1(_04605_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09968_ (.A1(_04602_),
    .A2(_02648_),
    .B(_04659_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09969_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_04605_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09970_ (.A1(_04658_),
    .A2(_04660_),
    .A3(_04661_),
    .A4(_04607_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09971_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_04603_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09972_ (.I(_04663_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09973_ (.A1(_04662_),
    .A2(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09974_ (.A1(_04655_),
    .A2(_04665_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09975_ (.A1(_04654_),
    .A2(_04666_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09976_ (.A1(_04649_),
    .A2(_04667_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09977_ (.A1(_04608_),
    .A2(_04620_),
    .B1(_04625_),
    .B2(_04643_),
    .C(_04668_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09978_ (.I(_04599_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09979_ (.A1(_04281_),
    .A2(_04670_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09980_ (.A1(_04601_),
    .A2(_04669_),
    .B(_04671_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09981_ (.I(_04660_),
    .Z(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09982_ (.I(_04629_),
    .Z(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09983_ (.I(_04598_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09984_ (.A1(_04672_),
    .A2(_04620_),
    .B1(_04625_),
    .B2(_04673_),
    .C(_04674_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09985_ (.A1(_02542_),
    .A2(_04601_),
    .B(_04675_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09986_ (.I(_03277_),
    .Z(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09987_ (.I(_04676_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09988_ (.A1(_02707_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09989_ (.A1(_04596_),
    .A2(\u_arbiter.i_wb_cpu_rdt[4] ),
    .B(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09990_ (.I(_03277_),
    .Z(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09991_ (.I(_04619_),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09992_ (.A1(_04680_),
    .A2(_04681_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09993_ (.I(_04682_),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09994_ (.I(_04653_),
    .Z(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09995_ (.A1(_04649_),
    .A2(_04684_),
    .A3(_04665_),
    .Z(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09996_ (.I(_04622_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09997_ (.I(_04655_),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09998_ (.A1(_04686_),
    .A2(_04687_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09999_ (.I(_04650_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10000_ (.I(_04627_),
    .Z(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10001_ (.I(_04663_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10002_ (.A1(_04655_),
    .A2(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10003_ (.A1(_04655_),
    .A2(_04690_),
    .B(_04692_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10004_ (.A1(_04612_),
    .A2(_04618_),
    .Z(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10005_ (.A1(_03277_),
    .A2(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10006_ (.A1(_04689_),
    .A2(_04693_),
    .B(_04695_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10007_ (.A1(_04685_),
    .A2(_04688_),
    .A3(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10008_ (.A1(_02557_),
    .A2(_04677_),
    .B1(_04679_),
    .B2(_04683_),
    .C(_04697_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10009_ (.I(_04680_),
    .Z(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10010_ (.I(_04698_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10011_ (.A1(_04609_),
    .A2(_04653_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10012_ (.I(_04700_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10013_ (.A1(_04616_),
    .A2(_04690_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10014_ (.I(_04634_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10015_ (.A1(_04703_),
    .A2(_04635_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10016_ (.I(_04640_),
    .Z(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10017_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_02706_),
    .Z(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10018_ (.A1(_04604_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10019_ (.A1(_03274_),
    .A2(\u_arbiter.i_wb_cpu_rdt[14] ),
    .B(_04707_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10020_ (.A1(_04708_),
    .A2(_04691_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10021_ (.A1(_04638_),
    .A2(_04705_),
    .B(_04706_),
    .C(_04709_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10022_ (.I(_04693_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10023_ (.A1(_04702_),
    .A2(_04704_),
    .B(_04710_),
    .C(_04711_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10024_ (.I(_04630_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10025_ (.I(_04713_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10026_ (.A1(_02708_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10027_ (.A1(_04596_),
    .A2(\u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_04715_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10028_ (.I(_04598_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10029_ (.A1(_04686_),
    .A2(_04714_),
    .B1(_04620_),
    .B2(_04716_),
    .C(_04717_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10030_ (.A1(_04701_),
    .A2(_04712_),
    .B(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10031_ (.A1(_02627_),
    .A2(_04699_),
    .B(_04719_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10032_ (.I(_04680_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10033_ (.I(_04656_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10034_ (.I(_04721_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10035_ (.A1(_02617_),
    .A2(_04720_),
    .B1(_04722_),
    .B2(_04683_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10036_ (.A1(_04667_),
    .A2(_04696_),
    .B(_04723_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10037_ (.I(_04648_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10038_ (.A1(_04625_),
    .A2(_04673_),
    .B(_04681_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10039_ (.I(_04708_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10040_ (.A1(_04726_),
    .A2(_04630_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10041_ (.A1(_04622_),
    .A2(_04623_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10042_ (.I(_04657_),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10043_ (.A1(_04721_),
    .A2(_04729_),
    .B(_04704_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10044_ (.A1(_04708_),
    .A2(_04630_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10045_ (.I(_04731_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10046_ (.I(_04706_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10047_ (.A1(_04607_),
    .A2(_04642_),
    .B1(_04732_),
    .B2(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10048_ (.A1(_04702_),
    .A2(_04730_),
    .B(_04734_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10049_ (.A1(_04625_),
    .A2(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10050_ (.A1(_04724_),
    .A2(_04725_),
    .B1(_04727_),
    .B2(_04728_),
    .C(_04736_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10051_ (.A1(_04720_),
    .A2(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10052_ (.A1(_02493_),
    .A2(_04699_),
    .B(_04738_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10053_ (.I(_04694_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10054_ (.I(_04739_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10055_ (.A1(_04740_),
    .A2(_04688_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10056_ (.A1(_02707_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10057_ (.A1(_03275_),
    .A2(\u_arbiter.i_wb_cpu_rdt[10] ),
    .B(_04742_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10058_ (.A1(_04708_),
    .A2(_04691_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10059_ (.A1(_04744_),
    .A2(_04706_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10060_ (.A1(_04743_),
    .A2(_04721_),
    .B(_04745_),
    .C(_04703_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10061_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_04602_),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10062_ (.I(_04747_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10063_ (.I(_04629_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10064_ (.A1(_04748_),
    .A2(_04749_),
    .B1(_04642_),
    .B2(_04660_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10065_ (.A1(_04746_),
    .A2(_04750_),
    .B(_04701_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10066_ (.A1(_04740_),
    .A2(_04733_),
    .B1(_04741_),
    .B2(_04751_),
    .C(_04676_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10067_ (.A1(_02491_),
    .A2(_04699_),
    .B(_04752_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10068_ (.I(_04726_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10069_ (.A1(_04658_),
    .A2(_04704_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10070_ (.A1(_04702_),
    .A2(_04754_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10071_ (.A1(_04748_),
    .A2(_04749_),
    .B1(_04642_),
    .B2(_04661_),
    .C(_04755_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10072_ (.A1(_04753_),
    .A2(_04612_),
    .B1(_04701_),
    .B2(_04756_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10073_ (.A1(_04720_),
    .A2(_04757_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10074_ (.A1(_02522_),
    .A2(_04699_),
    .B(_04758_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10075_ (.A1(_04598_),
    .A2(_04694_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10076_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_02709_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10077_ (.A1(_04649_),
    .A2(_04666_),
    .B1(_04631_),
    .B2(_04608_),
    .C(_04684_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10078_ (.I(_04692_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10079_ (.A1(_04607_),
    .A2(_04690_),
    .A3(_04762_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10080_ (.I(_04747_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10081_ (.A1(_04764_),
    .A2(_04643_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10082_ (.A1(_04650_),
    .A2(_04763_),
    .A3(_04765_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10083_ (.A1(_04607_),
    .A2(_04732_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10084_ (.A1(_04617_),
    .A2(_04767_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10085_ (.A1(_03278_),
    .A2(_04612_),
    .A3(_04766_),
    .A4(_04768_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10086_ (.A1(_04761_),
    .A2(_04769_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10087_ (.A1(_04759_),
    .A2(_04760_),
    .B(_04770_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10088_ (.A1(_02539_),
    .A2(_04699_),
    .B(_04771_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10089_ (.I(_04759_),
    .Z(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10090_ (.I(_02707_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10091_ (.I(_04773_),
    .Z(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10092_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .S(_04774_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10093_ (.I(_04617_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10094_ (.I(_04732_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10095_ (.A1(_04672_),
    .A2(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10096_ (.A1(_04764_),
    .A2(_04642_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10097_ (.A1(_04650_),
    .A2(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10098_ (.I(_04709_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10099_ (.A1(_04691_),
    .A2(_04706_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10100_ (.A1(_04753_),
    .A2(_04782_),
    .B(_04653_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10101_ (.A1(_04650_),
    .A2(_04781_),
    .B(_04783_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10102_ (.A1(_04684_),
    .A2(_04780_),
    .B1(_04784_),
    .B2(_04660_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10103_ (.A1(_04776_),
    .A2(_04778_),
    .B(_04785_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10104_ (.I(_04680_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10105_ (.A1(_04772_),
    .A2(_04775_),
    .B1(_04786_),
    .B2(_04787_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10106_ (.A1(_01448_),
    .A2(_04677_),
    .B(_04788_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10107_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_02708_),
    .Z(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10108_ (.A1(_04622_),
    .A2(_04652_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10109_ (.I(_04790_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10110_ (.A1(_04721_),
    .A2(_04713_),
    .B1(_04616_),
    .B2(_04789_),
    .C1(_04777_),
    .C2(_04661_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10111_ (.A1(_04648_),
    .A2(_04710_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10112_ (.A1(_04726_),
    .A2(_04793_),
    .A3(_04782_),
    .B(_04624_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10113_ (.A1(_04728_),
    .A2(_04794_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10114_ (.A1(_04700_),
    .A2(_04779_),
    .B(_04679_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10115_ (.A1(_04795_),
    .A2(_04796_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10116_ (.A1(_04791_),
    .A2(_04792_),
    .B(_04797_),
    .C(_04739_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10117_ (.A1(_04740_),
    .A2(_04789_),
    .B(_04798_),
    .C(_04698_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10118_ (.A1(_02499_),
    .A2(_04677_),
    .B(_04799_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10119_ (.I(_04151_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10120_ (.A1(_02890_),
    .A2(_04426_),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10121_ (.I(_04801_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10122_ (.I(_04801_),
    .Z(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10123_ (.A1(\u_cpu.rf_ram.memory[114][0] ),
    .A2(_04803_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10124_ (.A1(_04800_),
    .A2(_04802_),
    .B(_04804_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10125_ (.I(_04157_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10126_ (.A1(\u_cpu.rf_ram.memory[114][1] ),
    .A2(_04803_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10127_ (.A1(_04805_),
    .A2(_04802_),
    .B(_04806_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10128_ (.I(_04160_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10129_ (.I(_04801_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10130_ (.A1(\u_cpu.rf_ram.memory[114][2] ),
    .A2(_04808_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10131_ (.A1(_04807_),
    .A2(_04802_),
    .B(_04809_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10132_ (.I(_04164_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10133_ (.A1(\u_cpu.rf_ram.memory[114][3] ),
    .A2(_04808_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10134_ (.A1(_04810_),
    .A2(_04802_),
    .B(_04811_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10135_ (.I(_04167_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10136_ (.A1(\u_cpu.rf_ram.memory[114][4] ),
    .A2(_04808_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10137_ (.A1(_04812_),
    .A2(_04802_),
    .B(_04813_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10138_ (.I(_04170_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(\u_cpu.rf_ram.memory[114][5] ),
    .A2(_04808_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10140_ (.A1(_04814_),
    .A2(_04803_),
    .B(_04815_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10141_ (.I(_04173_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10142_ (.A1(\u_cpu.rf_ram.memory[114][6] ),
    .A2(_04808_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10143_ (.A1(_04816_),
    .A2(_04803_),
    .B(_04817_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10144_ (.I(_04176_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10145_ (.A1(\u_cpu.rf_ram.memory[114][7] ),
    .A2(_04801_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10146_ (.A1(_04818_),
    .A2(_04803_),
    .B(_04819_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10147_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .S(_02708_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10148_ (.A1(_04613_),
    .A2(_04691_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10149_ (.A1(_04690_),
    .A2(_04821_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10150_ (.I(_04822_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10151_ (.A1(_04748_),
    .A2(_04823_),
    .B(_04624_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10152_ (.A1(_04648_),
    .A2(_04726_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10153_ (.A1(_04634_),
    .A2(_04743_),
    .A3(_04764_),
    .A4(_04745_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10154_ (.A1(_04782_),
    .A2(_04825_),
    .B(_04826_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10155_ (.A1(_04823_),
    .A2(_04827_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10156_ (.A1(_04764_),
    .A2(_04641_),
    .B(_04709_),
    .C(_04733_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10157_ (.A1(_04716_),
    .A2(_04641_),
    .B(_04829_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10158_ (.I(_04637_),
    .Z(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10159_ (.A1(_04831_),
    .A2(_04629_),
    .B1(_04732_),
    .B2(_04729_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10160_ (.I(_04832_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10161_ (.A1(_04828_),
    .A2(_04830_),
    .A3(_04833_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10162_ (.I(_04831_),
    .Z(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10163_ (.A1(_04608_),
    .A2(_04781_),
    .B1(_04777_),
    .B2(_04835_),
    .C(_04653_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10164_ (.A1(_04824_),
    .A2(_04834_),
    .B1(_04836_),
    .B2(_04689_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10165_ (.A1(_04753_),
    .A2(_04729_),
    .B1(_04744_),
    .B2(_04820_),
    .C1(_04727_),
    .C2(_04835_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10166_ (.A1(_04776_),
    .A2(_04838_),
    .B(_04695_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10167_ (.A1(_04759_),
    .A2(_04820_),
    .B1(_04837_),
    .B2(_04839_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10168_ (.A1(_01457_),
    .A2(_04677_),
    .B(_04840_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10169_ (.A1(_04281_),
    .A2(_02627_),
    .A3(_01445_),
    .B(_02461_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10170_ (.A1(_04599_),
    .A2(_04841_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10171_ (.I(_04842_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10172_ (.A1(_04676_),
    .A2(_04841_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10173_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_04843_),
    .B1(_04844_),
    .B2(\u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10174_ (.A1(_04771_),
    .A2(_04845_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10175_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_04843_),
    .B1(_04844_),
    .B2(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10176_ (.A1(_04788_),
    .A2(_04846_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10177_ (.I(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10178_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_04841_),
    .B(_04674_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10179_ (.A1(_04847_),
    .A2(_04843_),
    .B1(_04848_),
    .B2(_04799_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10180_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .S(_02708_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10181_ (.I(_04790_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10182_ (.A1(_04702_),
    .A2(_04704_),
    .B(_04779_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10183_ (.I(_04794_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10184_ (.A1(_04729_),
    .A2(_04795_),
    .B1(_04851_),
    .B2(_04852_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10185_ (.A1(_04743_),
    .A2(_04713_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10186_ (.A1(_04687_),
    .A2(_04854_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10187_ (.A1(_04729_),
    .A2(_04821_),
    .B1(_04849_),
    .B2(_04664_),
    .C(_04790_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10188_ (.A1(_04850_),
    .A2(_04853_),
    .B1(_04855_),
    .B2(_04856_),
    .C(_04681_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10189_ (.A1(_04620_),
    .A2(_04849_),
    .B(_04857_),
    .C(_04600_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10190_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_04787_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10191_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_04843_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10192_ (.A1(_04843_),
    .A2(_04858_),
    .A3(_04859_),
    .B(_04860_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10193_ (.I(_04695_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10194_ (.I(_04703_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10195_ (.I(_04712_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10196_ (.A1(_04862_),
    .A2(_04673_),
    .B1(_04863_),
    .B2(_04722_),
    .C(_04780_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10197_ (.I(_04616_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10198_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_04773_),
    .Z(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10199_ (.A1(_04862_),
    .A2(_04714_),
    .B1(_04865_),
    .B2(_04866_),
    .C(_04791_),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10200_ (.A1(_04686_),
    .A2(_04722_),
    .B(_04684_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10201_ (.A1(_04861_),
    .A2(_04864_),
    .A3(_04867_),
    .A4(_04868_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10202_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_04842_),
    .B1(_04844_),
    .B2(\u_cpu.cpu.immdec.imm30_25[0] ),
    .C1(_04866_),
    .C2(_04772_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10203_ (.A1(_04869_),
    .A2(_04870_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10204_ (.A1(_04638_),
    .A2(_04705_),
    .A3(_04690_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10205_ (.A1(_04693_),
    .A2(_04871_),
    .B(_04608_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10206_ (.A1(_04748_),
    .A2(_04782_),
    .B(_04826_),
    .C(_04793_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10207_ (.A1(_04689_),
    .A2(_04872_),
    .A3(_04873_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10208_ (.A1(_04724_),
    .A2(_04686_),
    .B1(_04623_),
    .B2(_04688_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10209_ (.A1(_04874_),
    .A2(_04875_),
    .B(_04861_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10210_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .S(_04774_),
    .Z(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10211_ (.A1(_02614_),
    .A2(_02615_),
    .A3(_02463_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10212_ (.A1(_04281_),
    .A2(_04878_),
    .B(_02618_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10213_ (.A1(_03278_),
    .A2(_04879_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10214_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_04787_),
    .B1(_04682_),
    .B2(_04877_),
    .C(_04880_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10215_ (.A1(_03278_),
    .A2(_04879_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10216_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_04882_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10217_ (.A1(_04876_),
    .A2(_04881_),
    .B(_04883_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10218_ (.A1(_04717_),
    .A2(_04879_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10219_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_04882_),
    .B1(_04884_),
    .B2(\u_cpu.cpu.immdec.imm30_25[2] ),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10220_ (.A1(_04840_),
    .A2(_04885_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10221_ (.A1(_04672_),
    .A2(_04781_),
    .A3(_04871_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10222_ (.A1(_04722_),
    .A2(_04693_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10223_ (.A1(_04689_),
    .A2(_04873_),
    .A3(_04886_),
    .A4(_04887_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10224_ (.A1(_04644_),
    .A2(_04731_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10225_ (.A1(_04672_),
    .A2(_04781_),
    .B(_04684_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10226_ (.I(_04645_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10227_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_04773_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10228_ (.A1(_04891_),
    .A2(_04821_),
    .B1(_04892_),
    .B2(_04865_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10229_ (.A1(_04889_),
    .A2(_04890_),
    .B1(_04893_),
    .B2(_04776_),
    .C(_04695_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10230_ (.A1(_04888_),
    .A2(_04894_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10231_ (.A1(\u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_04882_),
    .B1(_04884_),
    .B2(\u_cpu.cpu.immdec.imm30_25[3] ),
    .C1(_04892_),
    .C2(_04772_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10232_ (.A1(_04895_),
    .A2(_04896_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10233_ (.I(_04636_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10234_ (.A1(_04897_),
    .A2(_04673_),
    .B1(_04777_),
    .B2(_04748_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10235_ (.A1(_04679_),
    .A2(_04641_),
    .B(_04829_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10236_ (.A1(_04828_),
    .A2(_04899_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10237_ (.A1(_04898_),
    .A2(_04900_),
    .B(_04824_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10238_ (.I(_04617_),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10239_ (.A1(_04897_),
    .A2(_04902_),
    .A3(_04821_),
    .Z(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10240_ (.A1(_04861_),
    .A2(_04901_),
    .A3(_04903_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10241_ (.A1(_04717_),
    .A2(_04879_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10242_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .S(_02709_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10243_ (.A1(\u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_04880_),
    .B1(_04905_),
    .B2(\u_cpu.cpu.immdec.imm30_25[4] ),
    .C1(_04906_),
    .C2(_04683_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10244_ (.A1(_04904_),
    .A2(_04907_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10245_ (.I(_04635_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10246_ (.A1(_04908_),
    .A2(_04673_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10247_ (.A1(_04724_),
    .A2(_04753_),
    .B(_04822_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10248_ (.A1(_04826_),
    .A2(_04910_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10249_ (.A1(_04909_),
    .A2(_04911_),
    .B(_04824_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10250_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .S(_04773_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10251_ (.A1(_04714_),
    .A2(_04913_),
    .B(_04854_),
    .C(_04902_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10252_ (.A1(_04687_),
    .A2(_04914_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10253_ (.A1(_04861_),
    .A2(_04912_),
    .A3(_04915_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _10254_ (.A1(\u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_04880_),
    .B1(_04905_),
    .B2(\u_cpu.cpu.immdec.imm30_25[5] ),
    .C1(_04913_),
    .C2(_04683_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10255_ (.A1(_04916_),
    .A2(_04917_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10256_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .S(_04774_),
    .Z(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10257_ (.A1(_04635_),
    .A2(_04724_),
    .B(_04703_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10258_ (.A1(_04862_),
    .A2(_04908_),
    .B1(_04754_),
    .B2(_04919_),
    .C(_04745_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10259_ (.A1(_04891_),
    .A2(_04749_),
    .B(_04910_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10260_ (.A1(_04920_),
    .A2(_04921_),
    .B(_04824_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10261_ (.A1(_04759_),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04698_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10262_ (.A1(\u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_04882_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10263_ (.I(\u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10264_ (.A1(_02614_),
    .A2(_04281_),
    .B(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10265_ (.A1(_02534_),
    .A2(_04926_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10266_ (.A1(_04925_),
    .A2(_04926_),
    .B(_04927_),
    .C(_02851_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10267_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_02851_),
    .B(_04884_),
    .C(_04928_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10268_ (.A1(_04923_),
    .A2(_04924_),
    .A3(_04929_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10269_ (.A1(_04831_),
    .A2(_04822_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10270_ (.A1(_04700_),
    .A2(_04930_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10271_ (.A1(_04637_),
    .A2(_04726_),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10272_ (.A1(_04831_),
    .A2(_04745_),
    .B1(_04932_),
    .B2(_04713_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10273_ (.A1(_04724_),
    .A2(_04762_),
    .B(_04933_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10274_ (.A1(_04646_),
    .A2(_04764_),
    .A3(_04666_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10275_ (.A1(_04831_),
    .A2(_04665_),
    .A3(_04692_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10276_ (.A1(_04623_),
    .A2(_04935_),
    .A3(_04936_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10277_ (.A1(_04931_),
    .A2(_04934_),
    .B1(_04937_),
    .B2(_04686_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10278_ (.A1(_04608_),
    .A2(_04714_),
    .B1(_04616_),
    .B2(_04835_),
    .C(_04850_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10279_ (.A1(_04938_),
    .A2(_04939_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10280_ (.A1(_04599_),
    .A2(_04681_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10281_ (.A1(_04835_),
    .A2(_04759_),
    .B1(_04940_),
    .B2(_04941_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10282_ (.A1(_02869_),
    .A2(_02534_),
    .B(_04674_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10283_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_02462_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10284_ (.A1(_04942_),
    .A2(_04943_),
    .B1(_04944_),
    .B2(_04601_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10285_ (.A1(_02614_),
    .A2(_02542_),
    .B(_02471_),
    .C(_02532_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10286_ (.A1(_02461_),
    .A2(_04945_),
    .B(_04680_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10287_ (.I(_04946_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10288_ (.I(_04947_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10289_ (.I(_04599_),
    .Z(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10290_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_04949_),
    .B(_04947_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10291_ (.A1(_04925_),
    .A2(_04948_),
    .B1(_04950_),
    .B2(_04771_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10292_ (.I(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10293_ (.I(_04946_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10294_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_04949_),
    .B(_04952_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10295_ (.A1(_04951_),
    .A2(_04948_),
    .B1(_04953_),
    .B2(_04738_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10296_ (.I(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10297_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_04949_),
    .B(_04952_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10298_ (.A1(_04954_),
    .A2(_04948_),
    .B1(_04955_),
    .B2(_04752_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10299_ (.I(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10300_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_04949_),
    .B(_04952_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10301_ (.A1(_04956_),
    .A2(_04948_),
    .B1(_04957_),
    .B2(_04758_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10302_ (.A1(_04747_),
    .A2(_04628_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10303_ (.A1(_04716_),
    .A2(_04710_),
    .B(_04958_),
    .C(_04823_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10304_ (.A1(_04931_),
    .A2(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10305_ (.A1(_04902_),
    .A2(_04727_),
    .A3(_04932_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10306_ (.A1(_04747_),
    .A2(_04662_),
    .A3(_04630_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10307_ (.A1(_04728_),
    .A2(_04655_),
    .A3(_04962_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10308_ (.A1(_04636_),
    .A2(_04822_),
    .B(_04624_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10309_ (.A1(_04713_),
    .A2(_04629_),
    .A3(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10310_ (.A1(_04963_),
    .A2(_04965_),
    .B(_04835_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10311_ (.A1(_04740_),
    .A2(_04960_),
    .A3(_04961_),
    .A4(_04966_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10312_ (.A1(_04664_),
    .A2(_04612_),
    .B(_04967_),
    .C(_04787_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10313_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_04670_),
    .B(_04947_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10314_ (.A1(_01439_),
    .A2(_04948_),
    .B1(_04968_),
    .B2(_04969_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10315_ (.I(_04952_),
    .Z(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10316_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .S(_04773_),
    .Z(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10317_ (.A1(_04865_),
    .A2(_04971_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10318_ (.A1(_04645_),
    .A2(_04687_),
    .B(_04790_),
    .C(_04821_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10319_ (.A1(_04733_),
    .A2(_04727_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10320_ (.A1(_04721_),
    .A2(_04641_),
    .B(_04709_),
    .C(_04733_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10321_ (.A1(_04645_),
    .A2(_04745_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10322_ (.A1(_04958_),
    .A2(_04822_),
    .A3(_04889_),
    .A4(_04976_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10323_ (.A1(_04705_),
    .A2(_04974_),
    .B1(_04975_),
    .B2(_04977_),
    .C(_04700_),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10324_ (.A1(_04705_),
    .A2(_04728_),
    .A3(_04962_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10325_ (.A1(_04790_),
    .A2(_04688_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10326_ (.A1(_04978_),
    .A2(_04979_),
    .A3(_04980_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10327_ (.A1(_04972_),
    .A2(_04973_),
    .B(_04681_),
    .C(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10328_ (.A1(_04620_),
    .A2(_04971_),
    .B(_04982_),
    .C(_04600_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10329_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_04698_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10330_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_04970_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10331_ (.A1(_04970_),
    .A2(_04983_),
    .A3(_04984_),
    .B(_04985_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10332_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_04970_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10333_ (.A1(_04596_),
    .A2(\u_arbiter.i_wb_cpu_rdt[17] ),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10334_ (.A1(_04596_),
    .A2(_02642_),
    .B(_04987_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10335_ (.A1(_04765_),
    .A2(_04823_),
    .B(_04964_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10336_ (.A1(_04963_),
    .A2(_04965_),
    .B(_04636_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10337_ (.A1(_04850_),
    .A2(_04990_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10338_ (.A1(_04989_),
    .A2(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10339_ (.A1(_04897_),
    .A2(_04687_),
    .B1(_04865_),
    .B2(_04988_),
    .C(_04850_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10340_ (.A1(_04992_),
    .A2(_04993_),
    .B(_04941_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10341_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_04676_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10342_ (.A1(_04952_),
    .A2(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10343_ (.A1(_04683_),
    .A2(_04988_),
    .B(_04994_),
    .C(_04996_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10344_ (.A1(_04986_),
    .A2(_04997_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10345_ (.A1(_04908_),
    .A2(_04963_),
    .B(_04617_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10346_ (.A1(_04749_),
    .A2(_04781_),
    .B(_04765_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10347_ (.A1(_04908_),
    .A2(_04823_),
    .B(_04999_),
    .C(_04625_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10348_ (.A1(_04753_),
    .A2(_04902_),
    .B1(_04998_),
    .B2(_05000_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10349_ (.A1(_04774_),
    .A2(\u_arbiter.i_wb_cpu_rdt[18] ),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10350_ (.A1(_02715_),
    .A2(_02646_),
    .B(_04739_),
    .C(_05002_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10351_ (.A1(_04600_),
    .A2(_05001_),
    .A3(_05003_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10352_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_04698_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10353_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_04947_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10354_ (.A1(_04970_),
    .A2(_05004_),
    .A3(_05005_),
    .B(_05006_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10355_ (.A1(_04703_),
    .A2(_04974_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10356_ (.A1(_04765_),
    .A2(_05007_),
    .B(_04701_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10357_ (.A1(_02709_),
    .A2(_02648_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10358_ (.A1(_04774_),
    .A2(\u_arbiter.i_wb_cpu_rdt[19] ),
    .B(_04619_),
    .C(_05009_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10359_ (.A1(_04676_),
    .A2(_05010_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10360_ (.A1(_04862_),
    .A2(_04963_),
    .B(_05008_),
    .C(_05011_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10361_ (.A1(_02616_),
    .A2(_01441_),
    .B(_04717_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10362_ (.A1(_02617_),
    .A2(_02534_),
    .B(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10363_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_04947_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10364_ (.A1(_04970_),
    .A2(_05012_),
    .A3(_05014_),
    .B(_05015_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10365_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .S(_02715_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10366_ (.A1(_04958_),
    .A2(_04911_),
    .B(_04824_),
    .C(_04717_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10367_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_04670_),
    .B1(_04772_),
    .B2(_05016_),
    .C(_05017_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10368_ (.I(_05018_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10369_ (.I(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10370_ (.A1(_04228_),
    .A2(_02874_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10371_ (.A1(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .A4(_05020_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10372_ (.A1(_05019_),
    .A2(_05020_),
    .B(_05021_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10373_ (.A1(_03067_),
    .A2(_03130_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10374_ (.I(_05022_),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10375_ (.I(_05022_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10376_ (.A1(\u_cpu.rf_ram.memory[32][0] ),
    .A2(_05024_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10377_ (.A1(_04800_),
    .A2(_05023_),
    .B(_05025_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10378_ (.A1(\u_cpu.rf_ram.memory[32][1] ),
    .A2(_05024_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10379_ (.A1(_04805_),
    .A2(_05023_),
    .B(_05026_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10380_ (.I(_05022_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10381_ (.A1(\u_cpu.rf_ram.memory[32][2] ),
    .A2(_05027_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10382_ (.A1(_04807_),
    .A2(_05023_),
    .B(_05028_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10383_ (.A1(\u_cpu.rf_ram.memory[32][3] ),
    .A2(_05027_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10384_ (.A1(_04810_),
    .A2(_05023_),
    .B(_05029_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(\u_cpu.rf_ram.memory[32][4] ),
    .A2(_05027_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10386_ (.A1(_04812_),
    .A2(_05023_),
    .B(_05030_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10387_ (.A1(\u_cpu.rf_ram.memory[32][5] ),
    .A2(_05027_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10388_ (.A1(_04814_),
    .A2(_05024_),
    .B(_05031_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10389_ (.A1(\u_cpu.rf_ram.memory[32][6] ),
    .A2(_05027_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10390_ (.A1(_04816_),
    .A2(_05024_),
    .B(_05032_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10391_ (.A1(\u_cpu.rf_ram.memory[32][7] ),
    .A2(_05022_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10392_ (.A1(_04818_),
    .A2(_05024_),
    .B(_05033_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10393_ (.A1(_03537_),
    .A2(_03231_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10394_ (.I(_05034_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10395_ (.I(_05034_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10396_ (.A1(\u_cpu.rf_ram.memory[31][0] ),
    .A2(_05036_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10397_ (.A1(_04800_),
    .A2(_05035_),
    .B(_05037_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10398_ (.A1(\u_cpu.rf_ram.memory[31][1] ),
    .A2(_05036_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10399_ (.A1(_04805_),
    .A2(_05035_),
    .B(_05038_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10400_ (.I(_05034_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10401_ (.A1(\u_cpu.rf_ram.memory[31][2] ),
    .A2(_05039_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10402_ (.A1(_04807_),
    .A2(_05035_),
    .B(_05040_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10403_ (.A1(\u_cpu.rf_ram.memory[31][3] ),
    .A2(_05039_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10404_ (.A1(_04810_),
    .A2(_05035_),
    .B(_05041_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10405_ (.A1(\u_cpu.rf_ram.memory[31][4] ),
    .A2(_05039_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10406_ (.A1(_04812_),
    .A2(_05035_),
    .B(_05042_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10407_ (.A1(\u_cpu.rf_ram.memory[31][5] ),
    .A2(_05039_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10408_ (.A1(_04814_),
    .A2(_05036_),
    .B(_05043_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10409_ (.A1(\u_cpu.rf_ram.memory[31][6] ),
    .A2(_05039_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10410_ (.A1(_04816_),
    .A2(_05036_),
    .B(_05044_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10411_ (.A1(\u_cpu.rf_ram.memory[31][7] ),
    .A2(_05034_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10412_ (.A1(_04818_),
    .A2(_05036_),
    .B(_05045_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10413_ (.A1(\u_cpu.cpu.alu.cmp_r ),
    .A2(_02869_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10414_ (.A1(_02869_),
    .A2(_04290_),
    .B(_05046_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10415_ (.I(_02530_),
    .Z(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10416_ (.I(_05047_),
    .Z(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10417_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_05048_),
    .Z(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10418_ (.I(_05049_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10419_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_05048_),
    .Z(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10420_ (.I(_05050_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10421_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_05048_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10422_ (.I(_05051_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10423_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_05048_),
    .Z(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10424_ (.I(_05052_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10425_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_05048_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10426_ (.I(_05053_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10427_ (.I(_05047_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10428_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_05054_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10429_ (.I(_05055_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10430_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_05054_),
    .Z(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10431_ (.I(_05056_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10432_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_05054_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10433_ (.I(_05057_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10434_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_05054_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10435_ (.I(_05058_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10436_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_05054_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10437_ (.I(_05059_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10438_ (.I(_05047_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10439_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_05060_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10440_ (.I(_05061_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10441_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_05060_),
    .Z(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10442_ (.I(_05062_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10443_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_05060_),
    .Z(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10444_ (.I(_05063_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10445_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_05060_),
    .Z(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10446_ (.I(_05064_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10447_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_05060_),
    .Z(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10448_ (.I(_05065_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10449_ (.I(_05047_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10450_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_05066_),
    .Z(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10451_ (.I(_05067_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10452_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_05066_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10453_ (.I(_05068_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10454_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_05066_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10455_ (.I(_05069_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10456_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_05066_),
    .Z(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10457_ (.I(_05070_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10458_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_05066_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10459_ (.I(_05071_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10460_ (.I(_05047_),
    .Z(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10461_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_05072_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10462_ (.I(_05073_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10463_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_05072_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10464_ (.I(_05074_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10465_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_05072_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10466_ (.I(_05075_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10467_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_05072_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10468_ (.I(_05076_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10469_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_05072_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10470_ (.I(_05077_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10471_ (.I(_02530_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10472_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_05078_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10473_ (.I(_05079_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10474_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_05078_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10475_ (.I(_05080_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10476_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .S(_05078_),
    .Z(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10477_ (.I(_05081_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10478_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .S(_05078_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10479_ (.I(_05082_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10480_ (.A1(_02856_),
    .A2(_02858_),
    .B(_02874_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10481_ (.A1(_02856_),
    .A2(_02858_),
    .B(_05083_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10482_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .A3(_02874_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10483_ (.A1(_05084_),
    .A2(_05085_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10484_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .I1(_05086_),
    .S(_05078_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10485_ (.I(_05087_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10486_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .B(_02501_),
    .C(_03281_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10487_ (.A1(_02862_),
    .A2(_03281_),
    .B(_05088_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10488_ (.A1(_02635_),
    .A2(_05089_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10489_ (.A1(_02644_),
    .A2(_05089_),
    .B(_05090_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10490_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_02874_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10491_ (.A1(_05084_),
    .A2(_05091_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10492_ (.I0(_02635_),
    .I1(_05092_),
    .S(_05089_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10493_ (.I(_05093_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10494_ (.A1(_03537_),
    .A2(_03083_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10495_ (.I(_05094_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10496_ (.I(_05094_),
    .Z(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10497_ (.A1(\u_cpu.rf_ram.memory[30][0] ),
    .A2(_05096_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10498_ (.A1(_04800_),
    .A2(_05095_),
    .B(_05097_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10499_ (.A1(\u_cpu.rf_ram.memory[30][1] ),
    .A2(_05096_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10500_ (.A1(_04805_),
    .A2(_05095_),
    .B(_05098_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10501_ (.I(_05094_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10502_ (.A1(\u_cpu.rf_ram.memory[30][2] ),
    .A2(_05099_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10503_ (.A1(_04807_),
    .A2(_05095_),
    .B(_05100_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10504_ (.A1(\u_cpu.rf_ram.memory[30][3] ),
    .A2(_05099_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10505_ (.A1(_04810_),
    .A2(_05095_),
    .B(_05101_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10506_ (.A1(\u_cpu.rf_ram.memory[30][4] ),
    .A2(_05099_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10507_ (.A1(_04812_),
    .A2(_05095_),
    .B(_05102_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10508_ (.A1(\u_cpu.rf_ram.memory[30][5] ),
    .A2(_05099_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10509_ (.A1(_04814_),
    .A2(_05096_),
    .B(_05103_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10510_ (.A1(\u_cpu.rf_ram.memory[30][6] ),
    .A2(_05099_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10511_ (.A1(_04816_),
    .A2(_05096_),
    .B(_05104_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10512_ (.A1(\u_cpu.rf_ram.memory[30][7] ),
    .A2(_05094_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10513_ (.A1(_04818_),
    .A2(_05096_),
    .B(_05105_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10514_ (.A1(_02461_),
    .A2(_02864_),
    .B(_03270_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10515_ (.I(_05106_),
    .Z(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10516_ (.I(_05107_),
    .Z(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10517_ (.A1(_03270_),
    .A2(_02865_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10518_ (.I(_05109_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10519_ (.I(_05110_),
    .Z(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10520_ (.A1(_02513_),
    .A2(_05108_),
    .B1(_05111_),
    .B2(_02699_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10521_ (.I(_05112_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10522_ (.A1(_02699_),
    .A2(_05108_),
    .B1(_05111_),
    .B2(_02710_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10523_ (.I(_05113_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10524_ (.A1(_02710_),
    .A2(_05108_),
    .B1(_05111_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10525_ (.I(_05114_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10526_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_05108_),
    .B1(_05111_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10527_ (.I(_05115_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10528_ (.I(_05107_),
    .Z(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10529_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_05116_),
    .B1(_05111_),
    .B2(_02725_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10530_ (.I(_05117_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10531_ (.I(_05110_),
    .Z(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10532_ (.A1(_02725_),
    .A2(_05116_),
    .B1(_05118_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10533_ (.I(_05119_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10534_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_05116_),
    .B1(_05118_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10535_ (.I(_05120_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10536_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_05116_),
    .B1(_05118_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10537_ (.I(_05121_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10538_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_05116_),
    .B1(_05118_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10539_ (.I(_05122_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10540_ (.I(_05106_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10541_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_05123_),
    .B1(_05118_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10542_ (.I(_05124_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10543_ (.I(_05110_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10544_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_05123_),
    .B1(_05125_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10545_ (.I(_05126_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10546_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_05123_),
    .B1(_05125_),
    .B2(_02758_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10547_ (.I(_05127_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10548_ (.A1(_02758_),
    .A2(_05123_),
    .B1(_05125_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10549_ (.I(_05128_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10550_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_05123_),
    .B1(_05125_),
    .B2(_02769_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10551_ (.I(_05129_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10552_ (.I(_05106_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10553_ (.A1(_02769_),
    .A2(_05130_),
    .B1(_05125_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10554_ (.I(_05131_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10555_ (.I(_05109_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10556_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_05130_),
    .B1(_05132_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10557_ (.I(_05133_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10558_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_05130_),
    .B1(_05132_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10559_ (.I(_05134_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10560_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_05130_),
    .B1(_05132_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10561_ (.I(_05135_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10562_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_05130_),
    .B1(_05132_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10563_ (.I(_05136_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10564_ (.I(_05106_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10565_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_05137_),
    .B1(_05132_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10566_ (.I(_05138_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10567_ (.I(_05109_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10568_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_05137_),
    .B1(_05139_),
    .B2(_02800_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10569_ (.I(_05140_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10570_ (.A1(_02800_),
    .A2(_05137_),
    .B1(_05139_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10571_ (.I(_05141_),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10572_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_05137_),
    .B1(_05139_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10573_ (.I(_05142_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10574_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_05137_),
    .B1(_05139_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10575_ (.I(_05143_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10576_ (.I(_05106_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10577_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_05144_),
    .B1(_05139_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10578_ (.I(_05145_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10579_ (.I(_05109_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10580_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_05144_),
    .B1(_05146_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10581_ (.I(_05147_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10582_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_05144_),
    .B1(_05146_),
    .B2(_02832_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10583_ (.I(_05148_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10584_ (.A1(_02832_),
    .A2(_05144_),
    .B1(_05146_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10585_ (.I(_05149_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10586_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_05144_),
    .B1(_05146_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10587_ (.I(_05150_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10588_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_05107_),
    .B1(_05146_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10589_ (.I(_05151_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10590_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_05107_),
    .B1(_05110_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10591_ (.I(_05152_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10592_ (.I0(_02577_),
    .I1(_02554_),
    .S(\u_cpu.cpu.ctrl.i_jump ),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10593_ (.A1(_02477_),
    .A2(_02548_),
    .B(_01454_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10594_ (.A1(_01454_),
    .A2(_05153_),
    .B(_05154_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10595_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_05107_),
    .B1(_05110_),
    .B2(_05155_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10596_ (.I(_05156_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10597_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_02897_),
    .A3(_03085_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10598_ (.I(_05157_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10599_ (.A1(_03131_),
    .A2(_05158_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10600_ (.I(_05159_),
    .Z(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10601_ (.I(_05159_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10602_ (.A1(\u_cpu.rf_ram.memory[109][0] ),
    .A2(_05161_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10603_ (.A1(_04800_),
    .A2(_05160_),
    .B(_05162_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10604_ (.A1(\u_cpu.rf_ram.memory[109][1] ),
    .A2(_05161_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10605_ (.A1(_04805_),
    .A2(_05160_),
    .B(_05163_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10606_ (.I(_05159_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10607_ (.A1(\u_cpu.rf_ram.memory[109][2] ),
    .A2(_05164_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10608_ (.A1(_04807_),
    .A2(_05160_),
    .B(_05165_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10609_ (.A1(\u_cpu.rf_ram.memory[109][3] ),
    .A2(_05164_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10610_ (.A1(_04810_),
    .A2(_05160_),
    .B(_05166_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10611_ (.A1(\u_cpu.rf_ram.memory[109][4] ),
    .A2(_05164_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10612_ (.A1(_04812_),
    .A2(_05160_),
    .B(_05167_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10613_ (.A1(\u_cpu.rf_ram.memory[109][5] ),
    .A2(_05164_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10614_ (.A1(_04814_),
    .A2(_05161_),
    .B(_05168_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10615_ (.A1(\u_cpu.rf_ram.memory[109][6] ),
    .A2(_05164_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10616_ (.A1(_04816_),
    .A2(_05161_),
    .B(_05169_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10617_ (.A1(\u_cpu.rf_ram.memory[109][7] ),
    .A2(_05159_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10618_ (.A1(_04818_),
    .A2(_05161_),
    .B(_05170_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10619_ (.A1(_03037_),
    .A2(_03480_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10620_ (.I(_05171_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10621_ (.I(_05171_),
    .Z(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10622_ (.A1(\u_cpu.rf_ram.memory[3][0] ),
    .A2(_05173_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10623_ (.A1(_04062_),
    .A2(_05172_),
    .B(_05174_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10624_ (.A1(\u_cpu.rf_ram.memory[3][1] ),
    .A2(_05173_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10625_ (.A1(_04068_),
    .A2(_05172_),
    .B(_05175_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10626_ (.I(_05171_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10627_ (.A1(\u_cpu.rf_ram.memory[3][2] ),
    .A2(_05176_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10628_ (.A1(_04070_),
    .A2(_05172_),
    .B(_05177_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10629_ (.A1(\u_cpu.rf_ram.memory[3][3] ),
    .A2(_05176_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10630_ (.A1(_04073_),
    .A2(_05172_),
    .B(_05178_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10631_ (.A1(\u_cpu.rf_ram.memory[3][4] ),
    .A2(_05176_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10632_ (.A1(_04075_),
    .A2(_05172_),
    .B(_05179_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10633_ (.A1(\u_cpu.rf_ram.memory[3][5] ),
    .A2(_05176_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10634_ (.A1(_04077_),
    .A2(_05173_),
    .B(_05180_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10635_ (.A1(\u_cpu.rf_ram.memory[3][6] ),
    .A2(_05176_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10636_ (.A1(_04079_),
    .A2(_05173_),
    .B(_05181_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10637_ (.A1(\u_cpu.rf_ram.memory[3][7] ),
    .A2(_05171_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10638_ (.A1(_04081_),
    .A2(_05173_),
    .B(_05182_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10639_ (.A1(_02891_),
    .A2(_03037_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10640_ (.I(_05183_),
    .Z(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10641_ (.I(_05183_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10642_ (.A1(\u_cpu.rf_ram.memory[2][0] ),
    .A2(_05185_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10643_ (.A1(_04062_),
    .A2(_05184_),
    .B(_05186_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10644_ (.A1(\u_cpu.rf_ram.memory[2][1] ),
    .A2(_05185_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10645_ (.A1(_04068_),
    .A2(_05184_),
    .B(_05187_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10646_ (.I(_05183_),
    .Z(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10647_ (.A1(\u_cpu.rf_ram.memory[2][2] ),
    .A2(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10648_ (.A1(_04070_),
    .A2(_05184_),
    .B(_05189_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10649_ (.A1(\u_cpu.rf_ram.memory[2][3] ),
    .A2(_05188_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10650_ (.A1(_04073_),
    .A2(_05184_),
    .B(_05190_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10651_ (.A1(\u_cpu.rf_ram.memory[2][4] ),
    .A2(_05188_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10652_ (.A1(_04075_),
    .A2(_05184_),
    .B(_05191_),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10653_ (.A1(\u_cpu.rf_ram.memory[2][5] ),
    .A2(_05188_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10654_ (.A1(_04077_),
    .A2(_05185_),
    .B(_05192_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10655_ (.A1(\u_cpu.rf_ram.memory[2][6] ),
    .A2(_05188_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10656_ (.A1(_04079_),
    .A2(_05185_),
    .B(_05193_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10657_ (.A1(\u_cpu.rf_ram.memory[2][7] ),
    .A2(_05183_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10658_ (.A1(_04081_),
    .A2(_05185_),
    .B(_05194_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10659_ (.I(_02905_),
    .Z(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10660_ (.I(_05195_),
    .Z(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10661_ (.A1(_04295_),
    .A2(_03132_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10662_ (.I(_05197_),
    .Z(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10663_ (.I(_05197_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10664_ (.A1(\u_cpu.rf_ram.memory[93][0] ),
    .A2(_05199_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10665_ (.A1(_05196_),
    .A2(_05198_),
    .B(_05200_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10666_ (.I(_02912_),
    .Z(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10667_ (.I(_05201_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10668_ (.A1(\u_cpu.rf_ram.memory[93][1] ),
    .A2(_05199_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10669_ (.A1(_05202_),
    .A2(_05198_),
    .B(_05203_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10670_ (.I(_02918_),
    .Z(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10671_ (.I(_05204_),
    .Z(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10672_ (.I(_05197_),
    .Z(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10673_ (.A1(\u_cpu.rf_ram.memory[93][2] ),
    .A2(_05206_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10674_ (.A1(_05205_),
    .A2(_05198_),
    .B(_05207_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10675_ (.I(_02925_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10676_ (.I(_05208_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10677_ (.A1(\u_cpu.rf_ram.memory[93][3] ),
    .A2(_05206_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10678_ (.A1(_05209_),
    .A2(_05198_),
    .B(_05210_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10679_ (.I(_02931_),
    .Z(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10680_ (.I(_05211_),
    .Z(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10681_ (.A1(\u_cpu.rf_ram.memory[93][4] ),
    .A2(_05206_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10682_ (.A1(_05212_),
    .A2(_05198_),
    .B(_05213_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10683_ (.I(_02937_),
    .Z(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10684_ (.I(_05214_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10685_ (.A1(\u_cpu.rf_ram.memory[93][5] ),
    .A2(_05206_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10686_ (.A1(_05215_),
    .A2(_05199_),
    .B(_05216_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10687_ (.I(_02943_),
    .Z(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10688_ (.I(_05217_),
    .Z(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10689_ (.A1(\u_cpu.rf_ram.memory[93][6] ),
    .A2(_05206_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10690_ (.A1(_05218_),
    .A2(_05199_),
    .B(_05219_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10691_ (.I(_02949_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10692_ (.I(_05220_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10693_ (.A1(\u_cpu.rf_ram.memory[93][7] ),
    .A2(_05197_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10694_ (.A1(_05221_),
    .A2(_05199_),
    .B(_05222_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10695_ (.A1(_02618_),
    .A2(_02873_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10696_ (.A1(_03278_),
    .A2(_05223_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10697_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_04674_),
    .B(_05224_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10698_ (.A1(_02467_),
    .A2(_05224_),
    .B1(_05225_),
    .B2(_04942_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10699_ (.A1(_04891_),
    .A2(_04654_),
    .A3(_04665_),
    .A4(_04762_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10700_ (.A1(_04645_),
    .A2(_04709_),
    .B1(_04732_),
    .B2(_04660_),
    .C(_04974_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10701_ (.A1(_04705_),
    .A2(_04974_),
    .B1(_04976_),
    .B2(_05227_),
    .C(_04700_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10702_ (.A1(_04776_),
    .A2(_05228_),
    .B(_04739_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10703_ (.A1(_04672_),
    .A2(_04714_),
    .B1(_04865_),
    .B2(_04891_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10704_ (.A1(_05226_),
    .A2(_05229_),
    .B1(_05230_),
    .B2(_04776_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10705_ (.A1(_04677_),
    .A2(_05231_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10706_ (.I(_05223_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10707_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_05233_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10708_ (.A1(_03084_),
    .A2(_05233_),
    .B(_05234_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10709_ (.A1(_04891_),
    .A2(_04772_),
    .B1(_05235_),
    .B2(_04670_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10710_ (.A1(_05232_),
    .A2(_05236_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10711_ (.A1(_04728_),
    .A2(_04666_),
    .B(_04739_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10712_ (.A1(_04897_),
    .A2(_05237_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10713_ (.A1(_04897_),
    .A2(_04711_),
    .A3(_04727_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10714_ (.A1(_04661_),
    .A2(_04777_),
    .B(_04974_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10715_ (.A1(_05239_),
    .A2(_05240_),
    .B(_04964_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10716_ (.A1(_04722_),
    .A2(_04902_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10717_ (.A1(_04679_),
    .A2(_04664_),
    .A3(_04791_),
    .B1(_04762_),
    .B2(_05242_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10718_ (.A1(_04674_),
    .A2(_05241_),
    .A3(_05243_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10719_ (.A1(_03084_),
    .A2(_05233_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10720_ (.A1(_02871_),
    .A2(_05233_),
    .B(_05245_),
    .C(_04787_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10721_ (.A1(_05238_),
    .A2(_05244_),
    .B(_05246_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10722_ (.A1(_02870_),
    .A2(_02618_),
    .A3(_02873_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10723_ (.A1(_02871_),
    .A2(_05233_),
    .B(_04949_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10724_ (.A1(_04623_),
    .A2(_04749_),
    .B(_04850_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10725_ (.A1(_05237_),
    .A2(_05249_),
    .B(_04908_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10726_ (.A1(_04664_),
    .A2(_04791_),
    .B1(_04701_),
    .B2(_04702_),
    .C(_05250_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10727_ (.A1(_04720_),
    .A2(_05251_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10728_ (.A1(_05247_),
    .A2(_05248_),
    .B(_05252_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10729_ (.A1(_04689_),
    .A2(_04631_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10730_ (.A1(_04782_),
    .A2(_05253_),
    .B(_04665_),
    .C(_04791_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10731_ (.A1(_04740_),
    .A2(_04762_),
    .A3(_05254_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10732_ (.A1(_04720_),
    .A2(_04862_),
    .A3(_05255_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10733_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_04670_),
    .B(_05224_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10734_ (.A1(_02894_),
    .A2(_05224_),
    .B1(_05256_),
    .B2(_05257_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(_02984_),
    .A2(_05158_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10736_ (.I(_05258_),
    .Z(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10737_ (.I(_05258_),
    .Z(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10738_ (.A1(\u_cpu.rf_ram.memory[97][0] ),
    .A2(_05260_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10739_ (.A1(_05196_),
    .A2(_05259_),
    .B(_05261_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10740_ (.A1(\u_cpu.rf_ram.memory[97][1] ),
    .A2(_05260_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10741_ (.A1(_05202_),
    .A2(_05259_),
    .B(_05262_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10742_ (.I(_05258_),
    .Z(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10743_ (.A1(\u_cpu.rf_ram.memory[97][2] ),
    .A2(_05263_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10744_ (.A1(_05205_),
    .A2(_05259_),
    .B(_05264_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10745_ (.A1(\u_cpu.rf_ram.memory[97][3] ),
    .A2(_05263_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10746_ (.A1(_05209_),
    .A2(_05259_),
    .B(_05265_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10747_ (.A1(\u_cpu.rf_ram.memory[97][4] ),
    .A2(_05263_),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10748_ (.A1(_05212_),
    .A2(_05259_),
    .B(_05266_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10749_ (.A1(\u_cpu.rf_ram.memory[97][5] ),
    .A2(_05263_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10750_ (.A1(_05215_),
    .A2(_05260_),
    .B(_05267_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10751_ (.A1(\u_cpu.rf_ram.memory[97][6] ),
    .A2(_05263_),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10752_ (.A1(_05218_),
    .A2(_05260_),
    .B(_05268_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10753_ (.A1(\u_cpu.rf_ram.memory[97][7] ),
    .A2(_05258_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10754_ (.A1(_05221_),
    .A2(_05260_),
    .B(_05269_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10755_ (.A1(_04295_),
    .A2(_03083_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10756_ (.I(_05270_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10757_ (.I(_05270_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10758_ (.A1(\u_cpu.rf_ram.memory[94][0] ),
    .A2(_05272_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10759_ (.A1(_05196_),
    .A2(_05271_),
    .B(_05273_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10760_ (.A1(\u_cpu.rf_ram.memory[94][1] ),
    .A2(_05272_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10761_ (.A1(_05202_),
    .A2(_05271_),
    .B(_05274_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10762_ (.I(_05270_),
    .Z(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10763_ (.A1(\u_cpu.rf_ram.memory[94][2] ),
    .A2(_05275_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10764_ (.A1(_05205_),
    .A2(_05271_),
    .B(_05276_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10765_ (.A1(\u_cpu.rf_ram.memory[94][3] ),
    .A2(_05275_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10766_ (.A1(_05209_),
    .A2(_05271_),
    .B(_05277_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10767_ (.A1(\u_cpu.rf_ram.memory[94][4] ),
    .A2(_05275_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10768_ (.A1(_05212_),
    .A2(_05271_),
    .B(_05278_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10769_ (.A1(\u_cpu.rf_ram.memory[94][5] ),
    .A2(_05275_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10770_ (.A1(_05215_),
    .A2(_05272_),
    .B(_05279_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10771_ (.A1(\u_cpu.rf_ram.memory[94][6] ),
    .A2(_05275_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10772_ (.A1(_05218_),
    .A2(_05272_),
    .B(_05280_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(\u_cpu.rf_ram.memory[94][7] ),
    .A2(_05270_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10774_ (.A1(_05221_),
    .A2(_05272_),
    .B(_05281_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10775_ (.A1(_04295_),
    .A2(_03231_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10776_ (.I(_05282_),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10777_ (.I(_05282_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10778_ (.A1(\u_cpu.rf_ram.memory[95][0] ),
    .A2(_05284_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10779_ (.A1(_05196_),
    .A2(_05283_),
    .B(_05285_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10780_ (.A1(\u_cpu.rf_ram.memory[95][1] ),
    .A2(_05284_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10781_ (.A1(_05202_),
    .A2(_05283_),
    .B(_05286_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10782_ (.I(_05282_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10783_ (.A1(\u_cpu.rf_ram.memory[95][2] ),
    .A2(_05287_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10784_ (.A1(_05205_),
    .A2(_05283_),
    .B(_05288_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10785_ (.A1(\u_cpu.rf_ram.memory[95][3] ),
    .A2(_05287_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10786_ (.A1(_05209_),
    .A2(_05283_),
    .B(_05289_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10787_ (.A1(\u_cpu.rf_ram.memory[95][4] ),
    .A2(_05287_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10788_ (.A1(_05212_),
    .A2(_05283_),
    .B(_05290_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10789_ (.A1(\u_cpu.rf_ram.memory[95][5] ),
    .A2(_05287_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10790_ (.A1(_05215_),
    .A2(_05284_),
    .B(_05291_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10791_ (.A1(\u_cpu.rf_ram.memory[95][6] ),
    .A2(_05287_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10792_ (.A1(_05218_),
    .A2(_05284_),
    .B(_05292_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10793_ (.A1(\u_cpu.rf_ram.memory[95][7] ),
    .A2(_05282_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10794_ (.A1(_05221_),
    .A2(_05284_),
    .B(_05293_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10795_ (.A1(_03067_),
    .A2(_05158_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10796_ (.I(_05294_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10797_ (.I(_05294_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10798_ (.A1(\u_cpu.rf_ram.memory[96][0] ),
    .A2(_05296_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10799_ (.A1(_05196_),
    .A2(_05295_),
    .B(_05297_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10800_ (.A1(\u_cpu.rf_ram.memory[96][1] ),
    .A2(_05296_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10801_ (.A1(_05202_),
    .A2(_05295_),
    .B(_05298_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10802_ (.I(_05294_),
    .Z(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10803_ (.A1(\u_cpu.rf_ram.memory[96][2] ),
    .A2(_05299_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10804_ (.A1(_05205_),
    .A2(_05295_),
    .B(_05300_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10805_ (.A1(\u_cpu.rf_ram.memory[96][3] ),
    .A2(_05299_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10806_ (.A1(_05209_),
    .A2(_05295_),
    .B(_05301_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10807_ (.A1(\u_cpu.rf_ram.memory[96][4] ),
    .A2(_05299_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10808_ (.A1(_05212_),
    .A2(_05295_),
    .B(_05302_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10809_ (.A1(\u_cpu.rf_ram.memory[96][5] ),
    .A2(_05299_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10810_ (.A1(_05215_),
    .A2(_05296_),
    .B(_05303_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10811_ (.A1(\u_cpu.rf_ram.memory[96][6] ),
    .A2(_05299_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10812_ (.A1(_05218_),
    .A2(_05296_),
    .B(_05304_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10813_ (.A1(\u_cpu.rf_ram.memory[96][7] ),
    .A2(_05294_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10814_ (.A1(_05221_),
    .A2(_05296_),
    .B(_05305_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10815_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_04601_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10816_ (.A1(_04923_),
    .A2(_05306_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10817_ (.A1(_02699_),
    .A2(_02632_),
    .A3(_02702_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10818_ (.A1(_02715_),
    .A2(_05307_),
    .Z(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10819_ (.A1(_03272_),
    .A2(_05308_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10820_ (.I(_05195_),
    .Z(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10821_ (.I(_02963_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10822_ (.A1(_05310_),
    .A2(_03153_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10823_ (.I(_05311_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10824_ (.I(_05311_),
    .Z(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10825_ (.A1(\u_cpu.rf_ram.memory[28][0] ),
    .A2(_05313_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10826_ (.A1(_05309_),
    .A2(_05312_),
    .B(_05314_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10827_ (.I(_05201_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10828_ (.A1(\u_cpu.rf_ram.memory[28][1] ),
    .A2(_05313_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10829_ (.A1(_05315_),
    .A2(_05312_),
    .B(_05316_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10830_ (.I(_05204_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10831_ (.I(_05311_),
    .Z(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10832_ (.A1(\u_cpu.rf_ram.memory[28][2] ),
    .A2(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10833_ (.A1(_05317_),
    .A2(_05312_),
    .B(_05319_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10834_ (.I(_05208_),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10835_ (.A1(\u_cpu.rf_ram.memory[28][3] ),
    .A2(_05318_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10836_ (.A1(_05320_),
    .A2(_05312_),
    .B(_05321_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10837_ (.I(_05211_),
    .Z(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10838_ (.A1(\u_cpu.rf_ram.memory[28][4] ),
    .A2(_05318_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10839_ (.A1(_05322_),
    .A2(_05312_),
    .B(_05323_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10840_ (.I(_05214_),
    .Z(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10841_ (.A1(\u_cpu.rf_ram.memory[28][5] ),
    .A2(_05318_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10842_ (.A1(_05324_),
    .A2(_05313_),
    .B(_05325_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10843_ (.I(_05217_),
    .Z(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10844_ (.A1(\u_cpu.rf_ram.memory[28][6] ),
    .A2(_05318_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10845_ (.A1(_05326_),
    .A2(_05313_),
    .B(_05327_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10846_ (.I(_05220_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10847_ (.A1(\u_cpu.rf_ram.memory[28][7] ),
    .A2(_05311_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10848_ (.A1(_05328_),
    .A2(_05313_),
    .B(_05329_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10849_ (.I(_03276_),
    .Z(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10850_ (.I(_05330_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10851_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_05331_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10852_ (.I(_05332_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10853_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_05331_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10854_ (.I(_05333_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10855_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_05331_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10856_ (.I(_05334_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10857_ (.I(_05330_),
    .Z(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10858_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_05335_),
    .Z(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10859_ (.I(_05336_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10860_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_05335_),
    .Z(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10861_ (.I(_05337_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10862_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_05335_),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10863_ (.I(_05338_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10864_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_05335_),
    .Z(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10865_ (.I(_05339_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10866_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_05335_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10867_ (.I(_05340_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10868_ (.I(_05330_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10869_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_05341_),
    .Z(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10870_ (.I(_05342_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10871_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_05341_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10872_ (.I(_05343_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10873_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_05341_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10874_ (.I(_05344_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10875_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_05331_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10876_ (.A1(_04632_),
    .A2(_05331_),
    .B(_05345_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10877_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_05341_),
    .Z(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10878_ (.I(_05346_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10879_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_05341_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10880_ (.I(_05347_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10881_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_05330_),
    .Z(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10882_ (.I(_05348_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10883_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_05330_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10884_ (.I(_05349_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10885_ (.A1(_02960_),
    .A2(_05158_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10886_ (.I(_05350_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10887_ (.I(_05350_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10888_ (.A1(\u_cpu.rf_ram.memory[101][0] ),
    .A2(_05352_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10889_ (.A1(_05309_),
    .A2(_05351_),
    .B(_05353_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10890_ (.A1(\u_cpu.rf_ram.memory[101][1] ),
    .A2(_05352_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10891_ (.A1(_05315_),
    .A2(_05351_),
    .B(_05354_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10892_ (.I(_05350_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10893_ (.A1(\u_cpu.rf_ram.memory[101][2] ),
    .A2(_05355_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10894_ (.A1(_05317_),
    .A2(_05351_),
    .B(_05356_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10895_ (.A1(\u_cpu.rf_ram.memory[101][3] ),
    .A2(_05355_),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10896_ (.A1(_05320_),
    .A2(_05351_),
    .B(_05357_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10897_ (.A1(\u_cpu.rf_ram.memory[101][4] ),
    .A2(_05355_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10898_ (.A1(_05322_),
    .A2(_05351_),
    .B(_05358_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10899_ (.A1(\u_cpu.rf_ram.memory[101][5] ),
    .A2(_05355_),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10900_ (.A1(_05324_),
    .A2(_05352_),
    .B(_05359_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10901_ (.A1(\u_cpu.rf_ram.memory[101][6] ),
    .A2(_05355_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10902_ (.A1(_05326_),
    .A2(_05352_),
    .B(_05360_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10903_ (.A1(\u_cpu.rf_ram.memory[101][7] ),
    .A2(_05350_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10904_ (.A1(_05328_),
    .A2(_05352_),
    .B(_05361_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10905_ (.A1(_03453_),
    .A2(_05158_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10906_ (.I(_05362_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10907_ (.I(_05362_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10908_ (.A1(\u_cpu.rf_ram.memory[102][0] ),
    .A2(_05364_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10909_ (.A1(_05309_),
    .A2(_05363_),
    .B(_05365_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10910_ (.A1(\u_cpu.rf_ram.memory[102][1] ),
    .A2(_05364_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10911_ (.A1(_05315_),
    .A2(_05363_),
    .B(_05366_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10912_ (.I(_05362_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10913_ (.A1(\u_cpu.rf_ram.memory[102][2] ),
    .A2(_05367_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10914_ (.A1(_05317_),
    .A2(_05363_),
    .B(_05368_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10915_ (.A1(\u_cpu.rf_ram.memory[102][3] ),
    .A2(_05367_),
    .ZN(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10916_ (.A1(_05320_),
    .A2(_05363_),
    .B(_05369_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10917_ (.A1(\u_cpu.rf_ram.memory[102][4] ),
    .A2(_05367_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10918_ (.A1(_05322_),
    .A2(_05363_),
    .B(_05370_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10919_ (.A1(\u_cpu.rf_ram.memory[102][5] ),
    .A2(_05367_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10920_ (.A1(_05324_),
    .A2(_05364_),
    .B(_05371_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10921_ (.A1(\u_cpu.rf_ram.memory[102][6] ),
    .A2(_05367_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10922_ (.A1(_05326_),
    .A2(_05364_),
    .B(_05372_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10923_ (.A1(\u_cpu.rf_ram.memory[102][7] ),
    .A2(_05362_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10924_ (.A1(_05328_),
    .A2(_05364_),
    .B(_05373_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10925_ (.I(_05157_),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10926_ (.A1(_03052_),
    .A2(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10927_ (.I(_05375_),
    .Z(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10928_ (.I(_05375_),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10929_ (.A1(\u_cpu.rf_ram.memory[103][0] ),
    .A2(_05377_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10930_ (.A1(_05309_),
    .A2(_05376_),
    .B(_05378_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10931_ (.A1(\u_cpu.rf_ram.memory[103][1] ),
    .A2(_05377_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10932_ (.A1(_05315_),
    .A2(_05376_),
    .B(_05379_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10933_ (.I(_05375_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10934_ (.A1(\u_cpu.rf_ram.memory[103][2] ),
    .A2(_05380_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10935_ (.A1(_05317_),
    .A2(_05376_),
    .B(_05381_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10936_ (.A1(\u_cpu.rf_ram.memory[103][3] ),
    .A2(_05380_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10937_ (.A1(_05320_),
    .A2(_05376_),
    .B(_05382_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10938_ (.A1(\u_cpu.rf_ram.memory[103][4] ),
    .A2(_05380_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10939_ (.A1(_05322_),
    .A2(_05376_),
    .B(_05383_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10940_ (.A1(\u_cpu.rf_ram.memory[103][5] ),
    .A2(_05380_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10941_ (.A1(_05324_),
    .A2(_05377_),
    .B(_05384_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10942_ (.A1(\u_cpu.rf_ram.memory[103][6] ),
    .A2(_05380_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10943_ (.A1(_05326_),
    .A2(_05377_),
    .B(_05385_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10944_ (.A1(\u_cpu.rf_ram.memory[103][7] ),
    .A2(_05375_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10945_ (.A1(_05328_),
    .A2(_05377_),
    .B(_05386_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10946_ (.A1(_03327_),
    .A2(_05374_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10947_ (.I(_05387_),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10948_ (.I(_05387_),
    .Z(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10949_ (.A1(\u_cpu.rf_ram.memory[104][0] ),
    .A2(_05389_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10950_ (.A1(_05309_),
    .A2(_05388_),
    .B(_05390_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10951_ (.A1(\u_cpu.rf_ram.memory[104][1] ),
    .A2(_05389_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10952_ (.A1(_05315_),
    .A2(_05388_),
    .B(_05391_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10953_ (.I(_05387_),
    .Z(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10954_ (.A1(\u_cpu.rf_ram.memory[104][2] ),
    .A2(_05392_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10955_ (.A1(_05317_),
    .A2(_05388_),
    .B(_05393_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10956_ (.A1(\u_cpu.rf_ram.memory[104][3] ),
    .A2(_05392_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10957_ (.A1(_05320_),
    .A2(_05388_),
    .B(_05394_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10958_ (.A1(\u_cpu.rf_ram.memory[104][4] ),
    .A2(_05392_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10959_ (.A1(_05322_),
    .A2(_05388_),
    .B(_05395_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10960_ (.A1(\u_cpu.rf_ram.memory[104][5] ),
    .A2(_05392_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10961_ (.A1(_05324_),
    .A2(_05389_),
    .B(_05396_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10962_ (.A1(\u_cpu.rf_ram.memory[104][6] ),
    .A2(_05392_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10963_ (.A1(_05326_),
    .A2(_05389_),
    .B(_05397_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10964_ (.A1(\u_cpu.rf_ram.memory[104][7] ),
    .A2(_05387_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10965_ (.A1(_05328_),
    .A2(_05389_),
    .B(_05398_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10966_ (.I(_05195_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10967_ (.A1(_03166_),
    .A2(_05374_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10968_ (.I(_05400_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10969_ (.I(_05400_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10970_ (.A1(\u_cpu.rf_ram.memory[99][0] ),
    .A2(_05402_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10971_ (.A1(_05399_),
    .A2(_05401_),
    .B(_05403_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10972_ (.I(_05201_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10973_ (.A1(\u_cpu.rf_ram.memory[99][1] ),
    .A2(_05402_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10974_ (.A1(_05404_),
    .A2(_05401_),
    .B(_05405_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10975_ (.I(_05204_),
    .Z(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10976_ (.I(_05400_),
    .Z(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10977_ (.A1(\u_cpu.rf_ram.memory[99][2] ),
    .A2(_05407_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10978_ (.A1(_05406_),
    .A2(_05401_),
    .B(_05408_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10979_ (.I(_05208_),
    .Z(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10980_ (.A1(\u_cpu.rf_ram.memory[99][3] ),
    .A2(_05407_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10981_ (.A1(_05409_),
    .A2(_05401_),
    .B(_05410_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10982_ (.I(_05211_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10983_ (.A1(\u_cpu.rf_ram.memory[99][4] ),
    .A2(_05407_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10984_ (.A1(_05411_),
    .A2(_05401_),
    .B(_05412_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10985_ (.I(_05214_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10986_ (.A1(\u_cpu.rf_ram.memory[99][5] ),
    .A2(_05407_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10987_ (.A1(_05413_),
    .A2(_05402_),
    .B(_05414_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10988_ (.I(_05217_),
    .Z(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10989_ (.A1(\u_cpu.rf_ram.memory[99][6] ),
    .A2(_05407_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10990_ (.A1(_05415_),
    .A2(_05402_),
    .B(_05416_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10991_ (.I(_05220_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10992_ (.A1(\u_cpu.rf_ram.memory[99][7] ),
    .A2(_05400_),
    .ZN(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10993_ (.A1(_05417_),
    .A2(_05402_),
    .B(_05418_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10994_ (.A1(_03086_),
    .A2(_03230_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10995_ (.I(_05419_),
    .Z(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10996_ (.I(_05419_),
    .Z(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10997_ (.A1(\u_cpu.rf_ram.memory[79][0] ),
    .A2(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10998_ (.A1(_05399_),
    .A2(_05420_),
    .B(_05422_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10999_ (.A1(\u_cpu.rf_ram.memory[79][1] ),
    .A2(_05421_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11000_ (.A1(_05404_),
    .A2(_05420_),
    .B(_05423_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11001_ (.I(_05419_),
    .Z(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11002_ (.A1(\u_cpu.rf_ram.memory[79][2] ),
    .A2(_05424_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11003_ (.A1(_05406_),
    .A2(_05420_),
    .B(_05425_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11004_ (.A1(\u_cpu.rf_ram.memory[79][3] ),
    .A2(_05424_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11005_ (.A1(_05409_),
    .A2(_05420_),
    .B(_05426_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11006_ (.A1(\u_cpu.rf_ram.memory[79][4] ),
    .A2(_05424_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11007_ (.A1(_05411_),
    .A2(_05420_),
    .B(_05427_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11008_ (.A1(\u_cpu.rf_ram.memory[79][5] ),
    .A2(_05424_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11009_ (.A1(_05413_),
    .A2(_05421_),
    .B(_05428_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11010_ (.A1(\u_cpu.rf_ram.memory[79][6] ),
    .A2(_05424_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11011_ (.A1(_05415_),
    .A2(_05421_),
    .B(_05429_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11012_ (.A1(\u_cpu.rf_ram.memory[79][7] ),
    .A2(_05419_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11013_ (.A1(_05417_),
    .A2(_05421_),
    .B(_05430_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11014_ (.A1(_03182_),
    .A2(_05374_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11015_ (.I(_05431_),
    .Z(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11016_ (.I(_05431_),
    .Z(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11017_ (.A1(\u_cpu.rf_ram.memory[105][0] ),
    .A2(_05433_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11018_ (.A1(_05399_),
    .A2(_05432_),
    .B(_05434_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11019_ (.A1(\u_cpu.rf_ram.memory[105][1] ),
    .A2(_05433_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11020_ (.A1(_05404_),
    .A2(_05432_),
    .B(_05435_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11021_ (.I(_05431_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11022_ (.A1(\u_cpu.rf_ram.memory[105][2] ),
    .A2(_05436_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11023_ (.A1(_05406_),
    .A2(_05432_),
    .B(_05437_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11024_ (.A1(\u_cpu.rf_ram.memory[105][3] ),
    .A2(_05436_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11025_ (.A1(_05409_),
    .A2(_05432_),
    .B(_05438_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11026_ (.A1(\u_cpu.rf_ram.memory[105][4] ),
    .A2(_05436_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11027_ (.A1(_05411_),
    .A2(_05432_),
    .B(_05439_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11028_ (.A1(\u_cpu.rf_ram.memory[105][5] ),
    .A2(_05436_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11029_ (.A1(_05413_),
    .A2(_05433_),
    .B(_05440_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11030_ (.A1(\u_cpu.rf_ram.memory[105][6] ),
    .A2(_05436_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11031_ (.A1(_05415_),
    .A2(_05433_),
    .B(_05441_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11032_ (.A1(\u_cpu.rf_ram.memory[105][7] ),
    .A2(_05431_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11033_ (.A1(_05417_),
    .A2(_05433_),
    .B(_05442_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11034_ (.A1(_03101_),
    .A2(_05374_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11035_ (.I(_05443_),
    .Z(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11036_ (.I(_05443_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11037_ (.A1(\u_cpu.rf_ram.memory[106][0] ),
    .A2(_05445_),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11038_ (.A1(_05399_),
    .A2(_05444_),
    .B(_05446_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11039_ (.A1(\u_cpu.rf_ram.memory[106][1] ),
    .A2(_05445_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11040_ (.A1(_05404_),
    .A2(_05444_),
    .B(_05447_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11041_ (.I(_05443_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11042_ (.A1(\u_cpu.rf_ram.memory[106][2] ),
    .A2(_05448_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11043_ (.A1(_05406_),
    .A2(_05444_),
    .B(_05449_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11044_ (.A1(\u_cpu.rf_ram.memory[106][3] ),
    .A2(_05448_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11045_ (.A1(_05409_),
    .A2(_05444_),
    .B(_05450_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11046_ (.A1(\u_cpu.rf_ram.memory[106][4] ),
    .A2(_05448_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11047_ (.A1(_05411_),
    .A2(_05444_),
    .B(_05451_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11048_ (.A1(\u_cpu.rf_ram.memory[106][5] ),
    .A2(_05448_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11049_ (.A1(_05413_),
    .A2(_05445_),
    .B(_05452_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11050_ (.A1(\u_cpu.rf_ram.memory[106][6] ),
    .A2(_05448_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11051_ (.A1(_05415_),
    .A2(_05445_),
    .B(_05453_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11052_ (.A1(\u_cpu.rf_ram.memory[106][7] ),
    .A2(_05443_),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11053_ (.A1(_05417_),
    .A2(_05445_),
    .B(_05454_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11054_ (.I(_05157_),
    .Z(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11055_ (.A1(_03196_),
    .A2(_05455_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11056_ (.I(_05456_),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11057_ (.I(_05456_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11058_ (.A1(\u_cpu.rf_ram.memory[107][0] ),
    .A2(_05458_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11059_ (.A1(_05399_),
    .A2(_05457_),
    .B(_05459_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11060_ (.A1(\u_cpu.rf_ram.memory[107][1] ),
    .A2(_05458_),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11061_ (.A1(_05404_),
    .A2(_05457_),
    .B(_05460_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11062_ (.I(_05456_),
    .Z(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11063_ (.A1(\u_cpu.rf_ram.memory[107][2] ),
    .A2(_05461_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11064_ (.A1(_05406_),
    .A2(_05457_),
    .B(_05462_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11065_ (.A1(\u_cpu.rf_ram.memory[107][3] ),
    .A2(_05461_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11066_ (.A1(_05409_),
    .A2(_05457_),
    .B(_05463_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11067_ (.A1(\u_cpu.rf_ram.memory[107][4] ),
    .A2(_05461_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11068_ (.A1(_05411_),
    .A2(_05457_),
    .B(_05464_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11069_ (.A1(\u_cpu.rf_ram.memory[107][5] ),
    .A2(_05461_),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11070_ (.A1(_05413_),
    .A2(_05458_),
    .B(_05465_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11071_ (.A1(\u_cpu.rf_ram.memory[107][6] ),
    .A2(_05461_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11072_ (.A1(_05415_),
    .A2(_05458_),
    .B(_05466_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11073_ (.A1(\u_cpu.rf_ram.memory[107][7] ),
    .A2(_05456_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11074_ (.A1(_05417_),
    .A2(_05458_),
    .B(_05467_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11075_ (.I(_05195_),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11076_ (.A1(_04295_),
    .A2(_03480_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11077_ (.I(_05469_),
    .Z(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11078_ (.I(_05469_),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11079_ (.A1(\u_cpu.rf_ram.memory[83][0] ),
    .A2(_05471_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11080_ (.A1(_05468_),
    .A2(_05470_),
    .B(_05472_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11081_ (.I(_05201_),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11082_ (.A1(\u_cpu.rf_ram.memory[83][1] ),
    .A2(_05471_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11083_ (.A1(_05473_),
    .A2(_05470_),
    .B(_05474_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11084_ (.I(_05204_),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11085_ (.I(_05469_),
    .Z(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11086_ (.A1(\u_cpu.rf_ram.memory[83][2] ),
    .A2(_05476_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11087_ (.A1(_05475_),
    .A2(_05470_),
    .B(_05477_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11088_ (.I(_05208_),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11089_ (.A1(\u_cpu.rf_ram.memory[83][3] ),
    .A2(_05476_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11090_ (.A1(_05478_),
    .A2(_05470_),
    .B(_05479_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11091_ (.I(_05211_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11092_ (.A1(\u_cpu.rf_ram.memory[83][4] ),
    .A2(_05476_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11093_ (.A1(_05480_),
    .A2(_05470_),
    .B(_05481_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11094_ (.I(_05214_),
    .Z(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11095_ (.A1(\u_cpu.rf_ram.memory[83][5] ),
    .A2(_05476_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11096_ (.A1(_05482_),
    .A2(_05471_),
    .B(_05483_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11097_ (.I(_05217_),
    .Z(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11098_ (.A1(\u_cpu.rf_ram.memory[83][6] ),
    .A2(_05476_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11099_ (.A1(_05484_),
    .A2(_05471_),
    .B(_05485_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11100_ (.I(_05220_),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11101_ (.A1(\u_cpu.rf_ram.memory[83][7] ),
    .A2(_05469_),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11102_ (.A1(_05486_),
    .A2(_05471_),
    .B(_05487_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11103_ (.A1(_03152_),
    .A2(_05455_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11104_ (.I(_05488_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11105_ (.I(_05488_),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11106_ (.A1(\u_cpu.rf_ram.memory[108][0] ),
    .A2(_05490_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11107_ (.A1(_05468_),
    .A2(_05489_),
    .B(_05491_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11108_ (.A1(\u_cpu.rf_ram.memory[108][1] ),
    .A2(_05490_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11109_ (.A1(_05473_),
    .A2(_05489_),
    .B(_05492_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11110_ (.I(_05488_),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11111_ (.A1(\u_cpu.rf_ram.memory[108][2] ),
    .A2(_05493_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11112_ (.A1(_05475_),
    .A2(_05489_),
    .B(_05494_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11113_ (.A1(\u_cpu.rf_ram.memory[108][3] ),
    .A2(_05493_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11114_ (.A1(_05478_),
    .A2(_05489_),
    .B(_05495_),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11115_ (.A1(\u_cpu.rf_ram.memory[108][4] ),
    .A2(_05493_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11116_ (.A1(_05480_),
    .A2(_05489_),
    .B(_05496_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11117_ (.A1(\u_cpu.rf_ram.memory[108][5] ),
    .A2(_05493_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11118_ (.A1(_05482_),
    .A2(_05490_),
    .B(_05497_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11119_ (.A1(\u_cpu.rf_ram.memory[108][6] ),
    .A2(_05493_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11120_ (.A1(_05484_),
    .A2(_05490_),
    .B(_05498_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11121_ (.A1(\u_cpu.rf_ram.memory[108][7] ),
    .A2(_05488_),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11122_ (.A1(_05486_),
    .A2(_05490_),
    .B(_05499_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11123_ (.A1(_02960_),
    .A2(_03395_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11124_ (.I(_05500_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11125_ (.I(_05500_),
    .Z(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11126_ (.A1(\u_cpu.rf_ram.memory[69][0] ),
    .A2(_05502_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11127_ (.A1(_05468_),
    .A2(_05501_),
    .B(_05503_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11128_ (.A1(\u_cpu.rf_ram.memory[69][1] ),
    .A2(_05502_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11129_ (.A1(_05473_),
    .A2(_05501_),
    .B(_05504_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11130_ (.I(_05500_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11131_ (.A1(\u_cpu.rf_ram.memory[69][2] ),
    .A2(_05505_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11132_ (.A1(_05475_),
    .A2(_05501_),
    .B(_05506_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11133_ (.A1(\u_cpu.rf_ram.memory[69][3] ),
    .A2(_05505_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11134_ (.A1(_05478_),
    .A2(_05501_),
    .B(_05507_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11135_ (.A1(\u_cpu.rf_ram.memory[69][4] ),
    .A2(_05505_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11136_ (.A1(_05480_),
    .A2(_05501_),
    .B(_05508_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11137_ (.A1(\u_cpu.rf_ram.memory[69][5] ),
    .A2(_05505_),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11138_ (.A1(_05482_),
    .A2(_05502_),
    .B(_05509_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11139_ (.A1(\u_cpu.rf_ram.memory[69][6] ),
    .A2(_05505_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11140_ (.A1(_05484_),
    .A2(_05502_),
    .B(_05510_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11141_ (.A1(\u_cpu.rf_ram.memory[69][7] ),
    .A2(_05500_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11142_ (.A1(_05486_),
    .A2(_05502_),
    .B(_05511_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11143_ (.I(_02898_),
    .Z(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11144_ (.A1(_05512_),
    .A2(_03013_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11145_ (.I(_05513_),
    .Z(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11146_ (.I(_05513_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11147_ (.A1(\u_cpu.rf_ram.memory[84][0] ),
    .A2(_05515_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11148_ (.A1(_05468_),
    .A2(_05514_),
    .B(_05516_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11149_ (.A1(\u_cpu.rf_ram.memory[84][1] ),
    .A2(_05515_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11150_ (.A1(_05473_),
    .A2(_05514_),
    .B(_05517_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11151_ (.I(_05513_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11152_ (.A1(\u_cpu.rf_ram.memory[84][2] ),
    .A2(_05518_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11153_ (.A1(_05475_),
    .A2(_05514_),
    .B(_05519_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11154_ (.A1(\u_cpu.rf_ram.memory[84][3] ),
    .A2(_05518_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11155_ (.A1(_05478_),
    .A2(_05514_),
    .B(_05520_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11156_ (.A1(\u_cpu.rf_ram.memory[84][4] ),
    .A2(_05518_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11157_ (.A1(_05480_),
    .A2(_05514_),
    .B(_05521_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11158_ (.A1(\u_cpu.rf_ram.memory[84][5] ),
    .A2(_05518_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11159_ (.A1(_05482_),
    .A2(_05515_),
    .B(_05522_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11160_ (.A1(\u_cpu.rf_ram.memory[84][6] ),
    .A2(_05518_),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11161_ (.A1(_05484_),
    .A2(_05515_),
    .B(_05523_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11162_ (.A1(\u_cpu.rf_ram.memory[84][7] ),
    .A2(_05513_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11163_ (.A1(_05486_),
    .A2(_05515_),
    .B(_05524_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11164_ (.A1(_03167_),
    .A2(_03197_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11165_ (.I(_05525_),
    .Z(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11166_ (.I(_05525_),
    .Z(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11167_ (.A1(\u_cpu.rf_ram.memory[59][0] ),
    .A2(_05527_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11168_ (.A1(_05468_),
    .A2(_05526_),
    .B(_05528_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11169_ (.A1(\u_cpu.rf_ram.memory[59][1] ),
    .A2(_05527_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11170_ (.A1(_05473_),
    .A2(_05526_),
    .B(_05529_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11171_ (.I(_05525_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11172_ (.A1(\u_cpu.rf_ram.memory[59][2] ),
    .A2(_05530_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11173_ (.A1(_05475_),
    .A2(_05526_),
    .B(_05531_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11174_ (.A1(\u_cpu.rf_ram.memory[59][3] ),
    .A2(_05530_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11175_ (.A1(_05478_),
    .A2(_05526_),
    .B(_05532_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11176_ (.A1(\u_cpu.rf_ram.memory[59][4] ),
    .A2(_05530_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11177_ (.A1(_05480_),
    .A2(_05526_),
    .B(_05533_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11178_ (.A1(\u_cpu.rf_ram.memory[59][5] ),
    .A2(_05530_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11179_ (.A1(_05482_),
    .A2(_05527_),
    .B(_05534_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11180_ (.A1(\u_cpu.rf_ram.memory[59][6] ),
    .A2(_05530_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11181_ (.A1(_05484_),
    .A2(_05527_),
    .B(_05535_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11182_ (.A1(\u_cpu.rf_ram.memory[59][7] ),
    .A2(_05525_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11183_ (.A1(_05486_),
    .A2(_05527_),
    .B(_05536_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11184_ (.A1(_03256_),
    .A2(_03102_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11185_ (.I(_05537_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11186_ (.I(_05538_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11187_ (.I(_05538_),
    .Z(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11188_ (.A1(\u_cpu.rf_ram.memory[10][0] ),
    .A2(_05540_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11189_ (.A1(_02954_),
    .A2(_05539_),
    .B(_05541_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11190_ (.A1(\u_cpu.rf_ram.memory[10][1] ),
    .A2(_05540_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11191_ (.A1(_02969_),
    .A2(_05539_),
    .B(_05542_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11192_ (.I(_05538_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11193_ (.A1(\u_cpu.rf_ram.memory[10][2] ),
    .A2(_05543_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11194_ (.A1(_02971_),
    .A2(_05539_),
    .B(_05544_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11195_ (.A1(\u_cpu.rf_ram.memory[10][3] ),
    .A2(_05543_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11196_ (.A1(_02974_),
    .A2(_05539_),
    .B(_05545_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11197_ (.A1(\u_cpu.rf_ram.memory[10][4] ),
    .A2(_05543_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11198_ (.A1(_02976_),
    .A2(_05539_),
    .B(_05546_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11199_ (.A1(\u_cpu.rf_ram.memory[10][5] ),
    .A2(_05543_),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11200_ (.A1(_02978_),
    .A2(_05540_),
    .B(_05547_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11201_ (.A1(\u_cpu.rf_ram.memory[10][6] ),
    .A2(_05543_),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11202_ (.A1(_02980_),
    .A2(_05540_),
    .B(_05548_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11203_ (.A1(\u_cpu.rf_ram.memory[10][7] ),
    .A2(_05538_),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11204_ (.A1(_02982_),
    .A2(_05540_),
    .B(_05549_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11205_ (.I(_05195_),
    .Z(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11206_ (.A1(_05512_),
    .A2(_02961_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11207_ (.I(_05551_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11208_ (.I(_05551_),
    .Z(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11209_ (.A1(\u_cpu.rf_ram.memory[85][0] ),
    .A2(_05553_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11210_ (.A1(_05550_),
    .A2(_05552_),
    .B(_05554_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11211_ (.I(_05201_),
    .Z(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11212_ (.A1(\u_cpu.rf_ram.memory[85][1] ),
    .A2(_05553_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11213_ (.A1(_05555_),
    .A2(_05552_),
    .B(_05556_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11214_ (.I(_05204_),
    .Z(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11215_ (.I(_05551_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11216_ (.A1(\u_cpu.rf_ram.memory[85][2] ),
    .A2(_05558_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11217_ (.A1(_05557_),
    .A2(_05552_),
    .B(_05559_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11218_ (.I(_05208_),
    .Z(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11219_ (.A1(\u_cpu.rf_ram.memory[85][3] ),
    .A2(_05558_),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11220_ (.A1(_05560_),
    .A2(_05552_),
    .B(_05561_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11221_ (.I(_05211_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11222_ (.A1(\u_cpu.rf_ram.memory[85][4] ),
    .A2(_05558_),
    .ZN(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11223_ (.A1(_05562_),
    .A2(_05552_),
    .B(_05563_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11224_ (.I(_05214_),
    .Z(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11225_ (.A1(\u_cpu.rf_ram.memory[85][5] ),
    .A2(_05558_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11226_ (.A1(_05564_),
    .A2(_05553_),
    .B(_05565_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11227_ (.I(_05217_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11228_ (.A1(\u_cpu.rf_ram.memory[85][6] ),
    .A2(_05558_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11229_ (.A1(_05566_),
    .A2(_05553_),
    .B(_05567_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11230_ (.I(_05220_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11231_ (.A1(\u_cpu.rf_ram.memory[85][7] ),
    .A2(_05551_),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11232_ (.A1(_05568_),
    .A2(_05553_),
    .B(_05569_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11233_ (.A1(_03082_),
    .A2(_05455_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11234_ (.I(_05570_),
    .Z(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11235_ (.I(_05570_),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11236_ (.A1(\u_cpu.rf_ram.memory[110][0] ),
    .A2(_05572_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11237_ (.A1(_05550_),
    .A2(_05571_),
    .B(_05573_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11238_ (.A1(\u_cpu.rf_ram.memory[110][1] ),
    .A2(_05572_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11239_ (.A1(_05555_),
    .A2(_05571_),
    .B(_05574_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11240_ (.I(_05570_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11241_ (.A1(\u_cpu.rf_ram.memory[110][2] ),
    .A2(_05575_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11242_ (.A1(_05557_),
    .A2(_05571_),
    .B(_05576_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11243_ (.A1(\u_cpu.rf_ram.memory[110][3] ),
    .A2(_05575_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11244_ (.A1(_05560_),
    .A2(_05571_),
    .B(_05577_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11245_ (.A1(\u_cpu.rf_ram.memory[110][4] ),
    .A2(_05575_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11246_ (.A1(_05562_),
    .A2(_05571_),
    .B(_05578_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11247_ (.A1(\u_cpu.rf_ram.memory[110][5] ),
    .A2(_05575_),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11248_ (.A1(_05564_),
    .A2(_05572_),
    .B(_05579_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11249_ (.A1(\u_cpu.rf_ram.memory[110][6] ),
    .A2(_05575_),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11250_ (.A1(_05566_),
    .A2(_05572_),
    .B(_05580_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11251_ (.A1(\u_cpu.rf_ram.memory[110][7] ),
    .A2(_05570_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11252_ (.A1(_05568_),
    .A2(_05572_),
    .B(_05581_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11253_ (.A1(_05512_),
    .A2(_03453_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11254_ (.I(_05582_),
    .Z(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11255_ (.I(_05582_),
    .Z(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11256_ (.A1(\u_cpu.rf_ram.memory[86][0] ),
    .A2(_05584_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11257_ (.A1(_05550_),
    .A2(_05583_),
    .B(_05585_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11258_ (.A1(\u_cpu.rf_ram.memory[86][1] ),
    .A2(_05584_),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11259_ (.A1(_05555_),
    .A2(_05583_),
    .B(_05586_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11260_ (.I(_05582_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11261_ (.A1(\u_cpu.rf_ram.memory[86][2] ),
    .A2(_05587_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11262_ (.A1(_05557_),
    .A2(_05583_),
    .B(_05588_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11263_ (.A1(\u_cpu.rf_ram.memory[86][3] ),
    .A2(_05587_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11264_ (.A1(_05560_),
    .A2(_05583_),
    .B(_05589_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11265_ (.A1(\u_cpu.rf_ram.memory[86][4] ),
    .A2(_05587_),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11266_ (.A1(_05562_),
    .A2(_05583_),
    .B(_05590_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11267_ (.A1(\u_cpu.rf_ram.memory[86][5] ),
    .A2(_05587_),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11268_ (.A1(_05564_),
    .A2(_05584_),
    .B(_05591_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11269_ (.A1(\u_cpu.rf_ram.memory[86][6] ),
    .A2(_05587_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11270_ (.A1(_05566_),
    .A2(_05584_),
    .B(_05592_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11271_ (.A1(\u_cpu.rf_ram.memory[86][7] ),
    .A2(_05582_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11272_ (.A1(_05568_),
    .A2(_05584_),
    .B(_05593_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11273_ (.A1(_03230_),
    .A2(_05455_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11274_ (.I(_05594_),
    .Z(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11275_ (.I(_05594_),
    .Z(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11276_ (.A1(\u_cpu.rf_ram.memory[111][0] ),
    .A2(_05596_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11277_ (.A1(_05550_),
    .A2(_05595_),
    .B(_05597_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11278_ (.A1(\u_cpu.rf_ram.memory[111][1] ),
    .A2(_05596_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11279_ (.A1(_05555_),
    .A2(_05595_),
    .B(_05598_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11280_ (.I(_05594_),
    .Z(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11281_ (.A1(\u_cpu.rf_ram.memory[111][2] ),
    .A2(_05599_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11282_ (.A1(_05557_),
    .A2(_05595_),
    .B(_05600_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11283_ (.A1(\u_cpu.rf_ram.memory[111][3] ),
    .A2(_05599_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11284_ (.A1(_05560_),
    .A2(_05595_),
    .B(_05601_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11285_ (.A1(\u_cpu.rf_ram.memory[111][4] ),
    .A2(_05599_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11286_ (.A1(_05562_),
    .A2(_05595_),
    .B(_05602_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11287_ (.A1(\u_cpu.rf_ram.memory[111][5] ),
    .A2(_05599_),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11288_ (.A1(_05564_),
    .A2(_05596_),
    .B(_05603_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11289_ (.A1(\u_cpu.rf_ram.memory[111][6] ),
    .A2(_05599_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11290_ (.A1(_05566_),
    .A2(_05596_),
    .B(_05604_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11291_ (.A1(\u_cpu.rf_ram.memory[111][7] ),
    .A2(_05594_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11292_ (.A1(_05568_),
    .A2(_05596_),
    .B(_05605_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11293_ (.A1(_05512_),
    .A2(_03053_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11294_ (.I(_05606_),
    .Z(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11295_ (.I(_05606_),
    .Z(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11296_ (.A1(\u_cpu.rf_ram.memory[87][0] ),
    .A2(_05608_),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11297_ (.A1(_05550_),
    .A2(_05607_),
    .B(_05609_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11298_ (.A1(\u_cpu.rf_ram.memory[87][1] ),
    .A2(_05608_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11299_ (.A1(_05555_),
    .A2(_05607_),
    .B(_05610_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11300_ (.I(_05606_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11301_ (.A1(\u_cpu.rf_ram.memory[87][2] ),
    .A2(_05611_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11302_ (.A1(_05557_),
    .A2(_05607_),
    .B(_05612_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11303_ (.A1(\u_cpu.rf_ram.memory[87][3] ),
    .A2(_05611_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11304_ (.A1(_05560_),
    .A2(_05607_),
    .B(_05613_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11305_ (.A1(\u_cpu.rf_ram.memory[87][4] ),
    .A2(_05611_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11306_ (.A1(_05562_),
    .A2(_05607_),
    .B(_05614_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11307_ (.A1(\u_cpu.rf_ram.memory[87][5] ),
    .A2(_05611_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11308_ (.A1(_05564_),
    .A2(_05608_),
    .B(_05615_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11309_ (.A1(\u_cpu.rf_ram.memory[87][6] ),
    .A2(_05611_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11310_ (.A1(_05566_),
    .A2(_05608_),
    .B(_05616_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11311_ (.A1(\u_cpu.rf_ram.memory[87][7] ),
    .A2(_05606_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11312_ (.A1(_05568_),
    .A2(_05608_),
    .B(_05617_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11313_ (.I(_02906_),
    .Z(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11314_ (.A1(_05512_),
    .A2(_03328_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11315_ (.I(_05619_),
    .Z(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11316_ (.I(_05619_),
    .Z(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11317_ (.A1(\u_cpu.rf_ram.memory[88][0] ),
    .A2(_05621_),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11318_ (.A1(_05618_),
    .A2(_05620_),
    .B(_05622_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11319_ (.I(_02913_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11320_ (.A1(\u_cpu.rf_ram.memory[88][1] ),
    .A2(_05621_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11321_ (.A1(_05623_),
    .A2(_05620_),
    .B(_05624_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11322_ (.I(_02919_),
    .Z(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11323_ (.I(_05619_),
    .Z(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11324_ (.A1(\u_cpu.rf_ram.memory[88][2] ),
    .A2(_05626_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11325_ (.A1(_05625_),
    .A2(_05620_),
    .B(_05627_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11326_ (.I(_02926_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11327_ (.A1(\u_cpu.rf_ram.memory[88][3] ),
    .A2(_05626_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11328_ (.A1(_05628_),
    .A2(_05620_),
    .B(_05629_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11329_ (.I(_02932_),
    .Z(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11330_ (.A1(\u_cpu.rf_ram.memory[88][4] ),
    .A2(_05626_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11331_ (.A1(_05630_),
    .A2(_05620_),
    .B(_05631_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11332_ (.I(_02938_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11333_ (.A1(\u_cpu.rf_ram.memory[88][5] ),
    .A2(_05626_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11334_ (.A1(_05632_),
    .A2(_05621_),
    .B(_05633_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11335_ (.I(_02944_),
    .Z(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11336_ (.A1(\u_cpu.rf_ram.memory[88][6] ),
    .A2(_05626_),
    .ZN(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11337_ (.A1(_05634_),
    .A2(_05621_),
    .B(_05635_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11338_ (.I(_02950_),
    .Z(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11339_ (.A1(\u_cpu.rf_ram.memory[88][7] ),
    .A2(_05619_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11340_ (.A1(_05636_),
    .A2(_05621_),
    .B(_05637_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11341_ (.A1(_04228_),
    .A2(_02515_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11342_ (.A1(_02462_),
    .A2(_02507_),
    .A3(_02501_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11343_ (.A1(_05638_),
    .A2(_05639_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11344_ (.I(_05640_),
    .Z(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11345_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11346_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01442_),
    .A3(_01460_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11347_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_05643_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11348_ (.A1(_03273_),
    .A2(_05642_),
    .B(_05644_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11349_ (.A1(_05641_),
    .A2(_05645_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11350_ (.A1(_02504_),
    .A2(_05641_),
    .B(_05646_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11351_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .ZN(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11352_ (.A1(_02616_),
    .A2(_02627_),
    .B1(_05647_),
    .B2(_03273_),
    .C(_05644_),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11353_ (.A1(_05641_),
    .A2(_05648_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11354_ (.A1(_05642_),
    .A2(_05641_),
    .B(_05649_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11355_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11356_ (.A1(_05650_),
    .A2(_02515_),
    .B(_01461_),
    .C(_02617_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11357_ (.I0(_05651_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .S(_05640_),
    .Z(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11358_ (.I(_05652_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11359_ (.A1(_02539_),
    .A2(_05643_),
    .B(_05640_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11360_ (.A1(_05650_),
    .A2(_05641_),
    .B1(_05653_),
    .B2(_02512_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11361_ (.A1(_01461_),
    .A2(_02512_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11362_ (.A1(_04228_),
    .A2(_02507_),
    .B(_02515_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11363_ (.I0(_05654_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .S(_05655_),
    .Z(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11364_ (.I(_05656_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11365_ (.I(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11366_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_05638_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11367_ (.A1(_05657_),
    .A2(_05638_),
    .B(_05658_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11368_ (.I(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .ZN(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11369_ (.A1(_01449_),
    .A2(_04236_),
    .A3(_04233_),
    .A4(_02499_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11370_ (.A1(_02502_),
    .A2(_04232_),
    .A3(_05660_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11371_ (.A1(_02511_),
    .A2(_05661_),
    .B(_04234_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11372_ (.A1(_05659_),
    .A2(_05661_),
    .B(_05662_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11373_ (.A1(_01480_),
    .A2(_02503_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11374_ (.A1(_05657_),
    .A2(_01480_),
    .B(_02515_),
    .C(_05663_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11375_ (.A1(_01480_),
    .A2(_02511_),
    .B(_05664_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11376_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_05638_),
    .A3(_05663_),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11377_ (.A1(_05665_),
    .A2(_05666_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11378_ (.A1(\u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_04601_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11379_ (.A1(_04861_),
    .A2(_05667_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11380_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_04242_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11381_ (.A1(_03271_),
    .A2(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A3(_05021_),
    .B(_05668_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11382_ (.A1(_05310_),
    .A2(_03196_),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11383_ (.I(_05669_),
    .Z(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11384_ (.I(_05669_),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11385_ (.A1(\u_cpu.rf_ram.memory[27][0] ),
    .A2(_05671_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11386_ (.A1(_05618_),
    .A2(_05670_),
    .B(_05672_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11387_ (.A1(\u_cpu.rf_ram.memory[27][1] ),
    .A2(_05671_),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11388_ (.A1(_05623_),
    .A2(_05670_),
    .B(_05673_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11389_ (.I(_05669_),
    .Z(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11390_ (.A1(\u_cpu.rf_ram.memory[27][2] ),
    .A2(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11391_ (.A1(_05625_),
    .A2(_05670_),
    .B(_05675_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11392_ (.A1(\u_cpu.rf_ram.memory[27][3] ),
    .A2(_05674_),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11393_ (.A1(_05628_),
    .A2(_05670_),
    .B(_05676_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11394_ (.A1(\u_cpu.rf_ram.memory[27][4] ),
    .A2(_05674_),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11395_ (.A1(_05630_),
    .A2(_05670_),
    .B(_05677_),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11396_ (.A1(\u_cpu.rf_ram.memory[27][5] ),
    .A2(_05674_),
    .ZN(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11397_ (.A1(_05632_),
    .A2(_05671_),
    .B(_05678_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11398_ (.A1(\u_cpu.rf_ram.memory[27][6] ),
    .A2(_05674_),
    .ZN(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11399_ (.A1(_05634_),
    .A2(_05671_),
    .B(_05679_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11400_ (.A1(\u_cpu.rf_ram.memory[27][7] ),
    .A2(_05669_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11401_ (.A1(_05636_),
    .A2(_05671_),
    .B(_05680_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11402_ (.A1(_05310_),
    .A2(_03102_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11403_ (.I(_05681_),
    .Z(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11404_ (.I(_05681_),
    .Z(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11405_ (.A1(\u_cpu.rf_ram.memory[26][0] ),
    .A2(_05683_),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11406_ (.A1(_05618_),
    .A2(_05682_),
    .B(_05684_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11407_ (.A1(\u_cpu.rf_ram.memory[26][1] ),
    .A2(_05683_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11408_ (.A1(_05623_),
    .A2(_05682_),
    .B(_05685_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11409_ (.I(_05681_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11410_ (.A1(\u_cpu.rf_ram.memory[26][2] ),
    .A2(_05686_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11411_ (.A1(_05625_),
    .A2(_05682_),
    .B(_05687_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11412_ (.A1(\u_cpu.rf_ram.memory[26][3] ),
    .A2(_05686_),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11413_ (.A1(_05628_),
    .A2(_05682_),
    .B(_05688_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11414_ (.A1(\u_cpu.rf_ram.memory[26][4] ),
    .A2(_05686_),
    .ZN(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11415_ (.A1(_05630_),
    .A2(_05682_),
    .B(_05689_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11416_ (.A1(\u_cpu.rf_ram.memory[26][5] ),
    .A2(_05686_),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11417_ (.A1(_05632_),
    .A2(_05683_),
    .B(_05690_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11418_ (.A1(\u_cpu.rf_ram.memory[26][6] ),
    .A2(_05686_),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11419_ (.A1(_05634_),
    .A2(_05683_),
    .B(_05691_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11420_ (.A1(\u_cpu.rf_ram.memory[26][7] ),
    .A2(_05681_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11421_ (.A1(_05636_),
    .A2(_05683_),
    .B(_05692_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11422_ (.A1(_05310_),
    .A2(_03183_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11423_ (.I(_05693_),
    .Z(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11424_ (.I(_05693_),
    .Z(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11425_ (.A1(\u_cpu.rf_ram.memory[25][0] ),
    .A2(_05695_),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11426_ (.A1(_05618_),
    .A2(_05694_),
    .B(_05696_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11427_ (.A1(\u_cpu.rf_ram.memory[25][1] ),
    .A2(_05695_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11428_ (.A1(_05623_),
    .A2(_05694_),
    .B(_05697_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11429_ (.I(_05693_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11430_ (.A1(\u_cpu.rf_ram.memory[25][2] ),
    .A2(_05698_),
    .ZN(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11431_ (.A1(_05625_),
    .A2(_05694_),
    .B(_05699_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11432_ (.A1(\u_cpu.rf_ram.memory[25][3] ),
    .A2(_05698_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11433_ (.A1(_05628_),
    .A2(_05694_),
    .B(_05700_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11434_ (.A1(\u_cpu.rf_ram.memory[25][4] ),
    .A2(_05698_),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11435_ (.A1(_05630_),
    .A2(_05694_),
    .B(_05701_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11436_ (.A1(\u_cpu.rf_ram.memory[25][5] ),
    .A2(_05698_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11437_ (.A1(_05632_),
    .A2(_05695_),
    .B(_05702_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11438_ (.A1(\u_cpu.rf_ram.memory[25][6] ),
    .A2(_05698_),
    .ZN(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11439_ (.A1(_05634_),
    .A2(_05695_),
    .B(_05703_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11440_ (.A1(\u_cpu.rf_ram.memory[25][7] ),
    .A2(_05693_),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11441_ (.A1(_05636_),
    .A2(_05695_),
    .B(_05704_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11442_ (.A1(_05310_),
    .A2(_03327_),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11443_ (.I(_05705_),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11444_ (.I(_05705_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11445_ (.A1(\u_cpu.rf_ram.memory[24][0] ),
    .A2(_05707_),
    .ZN(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11446_ (.A1(_05618_),
    .A2(_05706_),
    .B(_05708_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11447_ (.A1(\u_cpu.rf_ram.memory[24][1] ),
    .A2(_05707_),
    .ZN(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11448_ (.A1(_05623_),
    .A2(_05706_),
    .B(_05709_),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11449_ (.I(_05705_),
    .Z(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11450_ (.A1(\u_cpu.rf_ram.memory[24][2] ),
    .A2(_05710_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11451_ (.A1(_05625_),
    .A2(_05706_),
    .B(_05711_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11452_ (.A1(\u_cpu.rf_ram.memory[24][3] ),
    .A2(_05710_),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11453_ (.A1(_05628_),
    .A2(_05706_),
    .B(_05712_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11454_ (.A1(\u_cpu.rf_ram.memory[24][4] ),
    .A2(_05710_),
    .ZN(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11455_ (.A1(_05630_),
    .A2(_05706_),
    .B(_05713_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11456_ (.A1(\u_cpu.rf_ram.memory[24][5] ),
    .A2(_05710_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11457_ (.A1(_05632_),
    .A2(_05707_),
    .B(_05714_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11458_ (.A1(\u_cpu.rf_ram.memory[24][6] ),
    .A2(_05710_),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11459_ (.A1(_05634_),
    .A2(_05707_),
    .B(_05715_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11460_ (.A1(\u_cpu.rf_ram.memory[24][7] ),
    .A2(_05705_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11461_ (.A1(_05636_),
    .A2(_05707_),
    .B(_05716_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11462_ (.A1(_03050_),
    .A2(_03068_),
    .Z(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11463_ (.I(_05717_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11464_ (.I(_05717_),
    .Z(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11465_ (.A1(\u_cpu.rf_ram.memory[0][0] ),
    .A2(_05719_),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11466_ (.A1(_02954_),
    .A2(_05718_),
    .B(_05720_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11467_ (.A1(\u_cpu.rf_ram.memory[0][1] ),
    .A2(_05719_),
    .ZN(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11468_ (.A1(_02969_),
    .A2(_05718_),
    .B(_05721_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11469_ (.I(_05717_),
    .Z(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11470_ (.A1(\u_cpu.rf_ram.memory[0][2] ),
    .A2(_05722_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11471_ (.A1(_02971_),
    .A2(_05718_),
    .B(_05723_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11472_ (.A1(\u_cpu.rf_ram.memory[0][3] ),
    .A2(_05722_),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11473_ (.A1(_02974_),
    .A2(_05718_),
    .B(_05724_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11474_ (.A1(\u_cpu.rf_ram.memory[0][4] ),
    .A2(_05722_),
    .ZN(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11475_ (.A1(_02976_),
    .A2(_05718_),
    .B(_05725_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11476_ (.A1(\u_cpu.rf_ram.memory[0][5] ),
    .A2(_05722_),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11477_ (.A1(_02978_),
    .A2(_05719_),
    .B(_05726_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11478_ (.A1(\u_cpu.rf_ram.memory[0][6] ),
    .A2(_05722_),
    .ZN(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11479_ (.A1(_02980_),
    .A2(_05719_),
    .B(_05727_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11480_ (.A1(\u_cpu.rf_ram.memory[0][7] ),
    .A2(_05717_),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11481_ (.A1(_02982_),
    .A2(_05719_),
    .B(_05728_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11482_ (.A1(_02890_),
    .A2(_05455_),
    .ZN(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11483_ (.I(_05729_),
    .Z(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11484_ (.I(_05729_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11485_ (.A1(\u_cpu.rf_ram.memory[98][0] ),
    .A2(_05731_),
    .ZN(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11486_ (.A1(_03620_),
    .A2(_05730_),
    .B(_05732_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11487_ (.A1(\u_cpu.rf_ram.memory[98][1] ),
    .A2(_05731_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11488_ (.A1(_03627_),
    .A2(_05730_),
    .B(_05733_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11489_ (.I(_05729_),
    .Z(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11490_ (.A1(\u_cpu.rf_ram.memory[98][2] ),
    .A2(_05734_),
    .ZN(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11491_ (.A1(_03630_),
    .A2(_05730_),
    .B(_05735_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11492_ (.A1(\u_cpu.rf_ram.memory[98][3] ),
    .A2(_05734_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11493_ (.A1(_03634_),
    .A2(_05730_),
    .B(_05736_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11494_ (.A1(\u_cpu.rf_ram.memory[98][4] ),
    .A2(_05734_),
    .ZN(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11495_ (.A1(_03637_),
    .A2(_05730_),
    .B(_05737_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11496_ (.A1(\u_cpu.rf_ram.memory[98][5] ),
    .A2(_05734_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11497_ (.A1(_03640_),
    .A2(_05731_),
    .B(_05738_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11498_ (.A1(\u_cpu.rf_ram.memory[98][6] ),
    .A2(_05734_),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11499_ (.A1(_03643_),
    .A2(_05731_),
    .B(_05739_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11500_ (.A1(\u_cpu.rf_ram.memory[98][7] ),
    .A2(_05729_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11501_ (.A1(_03646_),
    .A2(_05731_),
    .B(_05740_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11502_ (.A1(_03012_),
    .A2(_05157_),
    .ZN(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11503_ (.I(_05741_),
    .Z(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11504_ (.I(_05741_),
    .Z(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11505_ (.A1(\u_cpu.rf_ram.memory[100][0] ),
    .A2(_05743_),
    .ZN(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11506_ (.A1(_03620_),
    .A2(_05742_),
    .B(_05744_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11507_ (.A1(\u_cpu.rf_ram.memory[100][1] ),
    .A2(_05743_),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11508_ (.A1(_03627_),
    .A2(_05742_),
    .B(_05745_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11509_ (.I(_05741_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11510_ (.A1(\u_cpu.rf_ram.memory[100][2] ),
    .A2(_05746_),
    .ZN(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11511_ (.A1(_03630_),
    .A2(_05742_),
    .B(_05747_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11512_ (.A1(\u_cpu.rf_ram.memory[100][3] ),
    .A2(_05746_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11513_ (.A1(_03634_),
    .A2(_05742_),
    .B(_05748_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11514_ (.A1(\u_cpu.rf_ram.memory[100][4] ),
    .A2(_05746_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11515_ (.A1(_03637_),
    .A2(_05742_),
    .B(_05749_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11516_ (.A1(\u_cpu.rf_ram.memory[100][5] ),
    .A2(_05746_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11517_ (.A1(_03640_),
    .A2(_05743_),
    .B(_05750_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11518_ (.A1(\u_cpu.rf_ram.memory[100][6] ),
    .A2(_05746_),
    .ZN(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11519_ (.A1(_03643_),
    .A2(_05743_),
    .B(_05751_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11520_ (.A1(\u_cpu.rf_ram.memory[100][7] ),
    .A2(_05741_),
    .ZN(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11521_ (.A1(_03646_),
    .A2(_05743_),
    .B(_05752_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11522_ (.A1(_02898_),
    .A2(_03182_),
    .ZN(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11523_ (.I(_05753_),
    .Z(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11524_ (.I(_05753_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11525_ (.A1(\u_cpu.rf_ram.memory[89][0] ),
    .A2(_05755_),
    .ZN(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11526_ (.A1(_03620_),
    .A2(_05754_),
    .B(_05756_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11527_ (.A1(\u_cpu.rf_ram.memory[89][1] ),
    .A2(_05755_),
    .ZN(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11528_ (.A1(_03627_),
    .A2(_05754_),
    .B(_05757_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11529_ (.I(_05753_),
    .Z(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11530_ (.A1(\u_cpu.rf_ram.memory[89][2] ),
    .A2(_05758_),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11531_ (.A1(_03630_),
    .A2(_05754_),
    .B(_05759_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11532_ (.A1(\u_cpu.rf_ram.memory[89][3] ),
    .A2(_05758_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11533_ (.A1(_03634_),
    .A2(_05754_),
    .B(_05760_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11534_ (.A1(\u_cpu.rf_ram.memory[89][4] ),
    .A2(_05758_),
    .ZN(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11535_ (.A1(_03637_),
    .A2(_05754_),
    .B(_05761_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11536_ (.A1(\u_cpu.rf_ram.memory[89][5] ),
    .A2(_05758_),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11537_ (.A1(_03640_),
    .A2(_05755_),
    .B(_05762_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11538_ (.A1(\u_cpu.rf_ram.memory[89][6] ),
    .A2(_05758_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11539_ (.A1(_03643_),
    .A2(_05755_),
    .B(_05763_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11540_ (.A1(\u_cpu.rf_ram.memory[89][7] ),
    .A2(_05753_),
    .ZN(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11541_ (.A1(_03646_),
    .A2(_05755_),
    .B(_05764_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11542_ (.A1(_02963_),
    .A2(_03053_),
    .ZN(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11543_ (.I(_05765_),
    .Z(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11544_ (.I(_05765_),
    .Z(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11545_ (.A1(\u_cpu.rf_ram.memory[23][0] ),
    .A2(_05767_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11546_ (.A1(_03620_),
    .A2(_05766_),
    .B(_05768_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11547_ (.A1(\u_cpu.rf_ram.memory[23][1] ),
    .A2(_05767_),
    .ZN(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11548_ (.A1(_03627_),
    .A2(_05766_),
    .B(_05769_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11549_ (.I(_05765_),
    .Z(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11550_ (.A1(\u_cpu.rf_ram.memory[23][2] ),
    .A2(_05770_),
    .ZN(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11551_ (.A1(_03630_),
    .A2(_05766_),
    .B(_05771_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11552_ (.A1(\u_cpu.rf_ram.memory[23][3] ),
    .A2(_05770_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11553_ (.A1(_03634_),
    .A2(_05766_),
    .B(_05772_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11554_ (.A1(\u_cpu.rf_ram.memory[23][4] ),
    .A2(_05770_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11555_ (.A1(_03637_),
    .A2(_05766_),
    .B(_05773_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11556_ (.A1(\u_cpu.rf_ram.memory[23][5] ),
    .A2(_05770_),
    .ZN(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11557_ (.A1(_03640_),
    .A2(_05767_),
    .B(_05774_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11558_ (.A1(\u_cpu.rf_ram.memory[23][6] ),
    .A2(_05770_),
    .ZN(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11559_ (.A1(_03643_),
    .A2(_05767_),
    .B(_05775_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11560_ (.A1(\u_cpu.rf_ram.memory[23][7] ),
    .A2(_05765_),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11561_ (.A1(_03646_),
    .A2(_05767_),
    .B(_05776_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11562_ (.A1(_04600_),
    .A2(_04241_),
    .ZN(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11563_ (.A1(\u_cpu.cpu.state.ibus_cyc ),
    .A2(_05777_),
    .ZN(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11564_ (.A1(_05108_),
    .A2(_05777_),
    .B(_05778_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11565_ (.A1(_02585_),
    .A2(_02587_),
    .A3(\u_cpu.rf_ram.rdata[7] ),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11566_ (.I(_05779_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11567_ (.A1(_02585_),
    .A2(\u_cpu.rf_ram.rdata[7] ),
    .A3(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11568_ (.I(_05780_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11569_ (.A1(_04234_),
    .A2(\u_cpu.rf_ram_if.rreq_r ),
    .Z(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11570_ (.I(_05781_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11571_ (.A1(_02885_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .Z(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11572_ (.A1(_03279_),
    .A2(_05782_),
    .ZN(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11573_ (.A1(_03294_),
    .A2(_05783_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11574_ (.D(_00096_),
    .CLK(net209),
    .Q(\u_cpu.rf_ram.memory[82][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11575_ (.D(_00097_),
    .CLK(net209),
    .Q(\u_cpu.rf_ram.memory[82][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11576_ (.D(_00098_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[82][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11577_ (.D(_00099_),
    .CLK(net209),
    .Q(\u_cpu.rf_ram.memory[82][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11578_ (.D(_00100_),
    .CLK(net213),
    .Q(\u_cpu.rf_ram.memory[82][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11579_ (.D(_00101_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[82][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11580_ (.D(_00102_),
    .CLK(net213),
    .Q(\u_cpu.rf_ram.memory[82][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11581_ (.D(_00103_),
    .CLK(net214),
    .Q(\u_cpu.rf_ram.memory[82][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11582_ (.D(_00104_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11583_ (.D(_00105_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11584_ (.D(_00106_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11585_ (.D(_00107_),
    .CLK(net411),
    .Q(\u_cpu.rf_ram.memory[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11586_ (.D(_00108_),
    .CLK(net411),
    .Q(\u_cpu.rf_ram.memory[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11587_ (.D(_00109_),
    .CLK(net411),
    .Q(\u_cpu.rf_ram.memory[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11588_ (.D(_00110_),
    .CLK(net411),
    .Q(\u_cpu.rf_ram.memory[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11589_ (.D(_00111_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11590_ (.D(_00112_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[81][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11591_ (.D(_00113_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[81][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11592_ (.D(_00114_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[81][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11593_ (.D(_00115_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[81][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11594_ (.D(_00116_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[81][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11595_ (.D(_00117_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[81][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11596_ (.D(_00118_),
    .CLK(net215),
    .Q(\u_cpu.rf_ram.memory[81][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11597_ (.D(_00119_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[81][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11598_ (.D(_00120_),
    .CLK(net414),
    .Q(\u_cpu.rf_ram.memory[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11599_ (.D(_00121_),
    .CLK(net414),
    .Q(\u_cpu.rf_ram.memory[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11600_ (.D(_00122_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11601_ (.D(_00123_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11602_ (.D(_00124_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11603_ (.D(_00125_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11604_ (.D(_00126_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11605_ (.D(_00127_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11606_ (.D(_00128_),
    .CLK(net379),
    .Q(\u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11607_ (.D(_00129_),
    .CLK(net379),
    .Q(\u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11608_ (.D(_00130_),
    .CLK(net381),
    .Q(\u_cpu.rf_ram.memory[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11609_ (.D(_00131_),
    .CLK(net381),
    .Q(\u_cpu.rf_ram.memory[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11610_ (.D(_00132_),
    .CLK(net381),
    .Q(\u_cpu.rf_ram.memory[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11611_ (.D(_00133_),
    .CLK(net374),
    .Q(\u_cpu.rf_ram.memory[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11612_ (.D(_00134_),
    .CLK(net381),
    .Q(\u_cpu.rf_ram.memory[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11613_ (.D(_00135_),
    .CLK(net382),
    .Q(\u_cpu.rf_ram.memory[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11614_ (.D(_00136_),
    .CLK(net441),
    .Q(\u_cpu.rf_ram.memory[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11615_ (.D(_00137_),
    .CLK(net442),
    .Q(\u_cpu.rf_ram.memory[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11616_ (.D(_00138_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11617_ (.D(_00139_),
    .CLK(net504),
    .Q(\u_cpu.rf_ram.memory[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11618_ (.D(_00140_),
    .CLK(net498),
    .Q(\u_cpu.rf_ram.memory[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11619_ (.D(_00141_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11620_ (.D(_00142_),
    .CLK(net437),
    .Q(\u_cpu.rf_ram.memory[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11621_ (.D(_00143_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11622_ (.D(_00144_),
    .CLK(net209),
    .Q(\u_cpu.rf_ram.memory[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11623_ (.D(_00145_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11624_ (.D(_00146_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11625_ (.D(_00147_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11626_ (.D(_00148_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11627_ (.D(_00149_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11628_ (.D(_00150_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11629_ (.D(_00151_),
    .CLK(net209),
    .Q(\u_cpu.rf_ram.memory[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11630_ (.D(_00152_),
    .CLK(net187),
    .Q(\u_cpu.rf_ram.memory[80][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11631_ (.D(_00153_),
    .CLK(net190),
    .Q(\u_cpu.rf_ram.memory[80][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11632_ (.D(_00154_),
    .CLK(net208),
    .Q(\u_cpu.rf_ram.memory[80][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11633_ (.D(_00155_),
    .CLK(net208),
    .Q(\u_cpu.rf_ram.memory[80][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11634_ (.D(_00156_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[80][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11635_ (.D(_00157_),
    .CLK(net208),
    .Q(\u_cpu.rf_ram.memory[80][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11636_ (.D(_00158_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[80][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11637_ (.D(_00159_),
    .CLK(net190),
    .Q(\u_cpu.rf_ram.memory[80][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11638_ (.D(_00160_),
    .CLK(net163),
    .Q(\u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11639_ (.D(_00161_),
    .CLK(net163),
    .Q(\u_cpu.rf_ram.memory[78][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11640_ (.D(_00162_),
    .CLK(net166),
    .Q(\u_cpu.rf_ram.memory[78][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11641_ (.D(_00163_),
    .CLK(net163),
    .Q(\u_cpu.rf_ram.memory[78][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11642_ (.D(_00164_),
    .CLK(net163),
    .Q(\u_cpu.rf_ram.memory[78][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11643_ (.D(_00165_),
    .CLK(net164),
    .Q(\u_cpu.rf_ram.memory[78][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11644_ (.D(_00166_),
    .CLK(net163),
    .Q(\u_cpu.rf_ram.memory[78][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11645_ (.D(_00167_),
    .CLK(net164),
    .Q(\u_cpu.rf_ram.memory[78][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11646_ (.D(_00168_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[42][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11647_ (.D(_00169_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[42][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11648_ (.D(_00170_),
    .CLK(net395),
    .Q(\u_cpu.rf_ram.memory[42][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11649_ (.D(_00171_),
    .CLK(net395),
    .Q(\u_cpu.rf_ram.memory[42][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11650_ (.D(_00172_),
    .CLK(net395),
    .Q(\u_cpu.rf_ram.memory[42][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11651_ (.D(_00173_),
    .CLK(net389),
    .Q(\u_cpu.rf_ram.memory[42][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11652_ (.D(_00174_),
    .CLK(net389),
    .Q(\u_cpu.rf_ram.memory[42][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11653_ (.D(_00175_),
    .CLK(net389),
    .Q(\u_cpu.rf_ram.memory[42][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11654_ (.D(_00176_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11655_ (.D(_00177_),
    .CLK(net405),
    .Q(\u_cpu.rf_ram.memory[46][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11656_ (.D(_00178_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11657_ (.D(_00179_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[46][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11658_ (.D(_00180_),
    .CLK(net404),
    .Q(\u_cpu.rf_ram.memory[46][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11659_ (.D(_00181_),
    .CLK(net405),
    .Q(\u_cpu.rf_ram.memory[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11660_ (.D(_00182_),
    .CLK(net405),
    .Q(\u_cpu.rf_ram.memory[46][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11661_ (.D(_00183_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[46][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11662_ (.D(_00184_),
    .CLK(net463),
    .Q(\u_cpu.rf_ram.memory[45][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11663_ (.D(_00185_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[45][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11664_ (.D(_00186_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[45][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11665_ (.D(_00187_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[45][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11666_ (.D(_00188_),
    .CLK(net462),
    .Q(\u_cpu.rf_ram.memory[45][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11667_ (.D(_00189_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[45][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11668_ (.D(_00190_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[45][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11669_ (.D(_00191_),
    .CLK(net463),
    .Q(\u_cpu.rf_ram.memory[45][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11670_ (.D(_00192_),
    .CLK(net464),
    .Q(\u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11671_ (.D(_00193_),
    .CLK(net466),
    .Q(\u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11672_ (.D(_00194_),
    .CLK(net466),
    .Q(\u_cpu.rf_ram.memory[44][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11673_ (.D(_00195_),
    .CLK(net466),
    .Q(\u_cpu.rf_ram.memory[44][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11674_ (.D(_00196_),
    .CLK(net467),
    .Q(\u_cpu.rf_ram.memory[44][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11675_ (.D(_00197_),
    .CLK(net466),
    .Q(\u_cpu.rf_ram.memory[44][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11676_ (.D(_00198_),
    .CLK(net466),
    .Q(\u_cpu.rf_ram.memory[44][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11677_ (.D(_00199_),
    .CLK(net464),
    .Q(\u_cpu.rf_ram.memory[44][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11678_ (.D(_00200_),
    .CLK(net391),
    .Q(\u_cpu.rf_ram.memory[51][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11679_ (.D(_00201_),
    .CLK(net391),
    .Q(\u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11680_ (.D(_00202_),
    .CLK(net391),
    .Q(\u_cpu.rf_ram.memory[51][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11681_ (.D(_00203_),
    .CLK(net389),
    .Q(\u_cpu.rf_ram.memory[51][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11682_ (.D(_00204_),
    .CLK(net389),
    .Q(\u_cpu.rf_ram.memory[51][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11683_ (.D(_00205_),
    .CLK(net391),
    .Q(\u_cpu.rf_ram.memory[51][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11684_ (.D(_00206_),
    .CLK(net374),
    .Q(\u_cpu.rf_ram.memory[51][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00207_),
    .CLK(net374),
    .Q(\u_cpu.rf_ram.memory[51][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00208_),
    .CLK(net464),
    .Q(\u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00209_),
    .CLK(net464),
    .Q(\u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00210_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00211_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00212_),
    .CLK(net457),
    .Q(\u_cpu.rf_ram.memory[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00213_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00214_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00215_),
    .CLK(net457),
    .Q(\u_cpu.rf_ram.memory[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00216_),
    .CLK(net402),
    .Q(\u_cpu.rf_ram.memory[43][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00217_),
    .CLK(net402),
    .Q(\u_cpu.rf_ram.memory[43][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00218_),
    .CLK(net452),
    .Q(\u_cpu.rf_ram.memory[43][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11697_ (.D(_00219_),
    .CLK(net452),
    .Q(\u_cpu.rf_ram.memory[43][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00220_),
    .CLK(net453),
    .Q(\u_cpu.rf_ram.memory[43][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00221_),
    .CLK(net390),
    .Q(\u_cpu.rf_ram.memory[43][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00222_),
    .CLK(net390),
    .Q(\u_cpu.rf_ram.memory[43][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00223_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[43][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00224_),
    .CLK(net387),
    .Q(\u_cpu.rf_ram.memory[48][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00225_),
    .CLK(net387),
    .Q(\u_cpu.rf_ram.memory[48][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00226_),
    .CLK(net296),
    .Q(\u_cpu.rf_ram.memory[48][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00227_),
    .CLK(net393),
    .Q(\u_cpu.rf_ram.memory[48][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00228_),
    .CLK(net296),
    .Q(\u_cpu.rf_ram.memory[48][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00229_),
    .CLK(net388),
    .Q(\u_cpu.rf_ram.memory[48][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00230_),
    .CLK(net388),
    .Q(\u_cpu.rf_ram.memory[48][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00231_),
    .CLK(net374),
    .Q(\u_cpu.rf_ram.memory[48][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00232_),
    .CLK(net463),
    .Q(\u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00233_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[47][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00234_),
    .CLK(net404),
    .Q(\u_cpu.rf_ram.memory[47][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00235_),
    .CLK(net462),
    .Q(\u_cpu.rf_ram.memory[47][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00236_),
    .CLK(net462),
    .Q(\u_cpu.rf_ram.memory[47][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11715_ (.D(_00237_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00238_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[47][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00239_),
    .CLK(net402),
    .Q(\u_cpu.rf_ram.memory[47][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00240_),
    .CLK(net387),
    .Q(\u_cpu.rf_ram.memory[50][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00241_),
    .CLK(net387),
    .Q(\u_cpu.rf_ram.memory[50][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00242_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.memory[50][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00243_),
    .CLK(net387),
    .Q(\u_cpu.rf_ram.memory[50][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00244_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.memory[50][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00245_),
    .CLK(net375),
    .Q(\u_cpu.rf_ram.memory[50][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11724_ (.D(_00246_),
    .CLK(net375),
    .Q(\u_cpu.rf_ram.memory[50][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00247_),
    .CLK(net376),
    .Q(\u_cpu.rf_ram.memory[50][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00248_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00249_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00250_),
    .CLK(net218),
    .Q(\u_cpu.rf_ram.memory[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00251_),
    .CLK(net219),
    .Q(\u_cpu.rf_ram.memory[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00252_),
    .CLK(net219),
    .Q(\u_cpu.rf_ram.memory[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00253_),
    .CLK(net218),
    .Q(\u_cpu.rf_ram.memory[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00254_),
    .CLK(net218),
    .Q(\u_cpu.rf_ram.memory[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00255_),
    .CLK(net213),
    .Q(\u_cpu.rf_ram.memory[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00256_),
    .CLK(net316),
    .Q(\u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00257_),
    .CLK(net285),
    .Q(\u_cpu.rf_ram_if.rcnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00258_),
    .CLK(net337),
    .Q(\u_cpu.rf_ram_if.rcnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00259_),
    .CLK(net288),
    .Q(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00260_),
    .CLK(net288),
    .Q(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00261_),
    .CLK(net433),
    .Q(\u_cpu.rf_ram.memory[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00262_),
    .CLK(net433),
    .Q(\u_cpu.rf_ram.memory[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00263_),
    .CLK(net435),
    .Q(\u_cpu.rf_ram.memory[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00264_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00265_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00266_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00267_),
    .CLK(net431),
    .Q(\u_cpu.rf_ram.memory[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00268_),
    .CLK(net431),
    .Q(\u_cpu.rf_ram.memory[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00269_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00270_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00271_),
    .CLK(net429),
    .Q(\u_cpu.rf_ram.memory[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00272_),
    .CLK(net429),
    .Q(\u_cpu.rf_ram.memory[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00273_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00274_),
    .CLK(net429),
    .Q(\u_cpu.rf_ram.memory[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00275_),
    .CLK(net429),
    .Q(\u_cpu.rf_ram.memory[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00276_),
    .CLK(net429),
    .Q(\u_cpu.rf_ram.memory[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00277_),
    .CLK(net393),
    .Q(\u_cpu.rf_ram.memory[40][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00278_),
    .CLK(net393),
    .Q(\u_cpu.rf_ram.memory[40][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00279_),
    .CLK(net452),
    .Q(\u_cpu.rf_ram.memory[40][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00280_),
    .CLK(net453),
    .Q(\u_cpu.rf_ram.memory[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00281_),
    .CLK(net453),
    .Q(\u_cpu.rf_ram.memory[40][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00282_),
    .CLK(net396),
    .Q(\u_cpu.rf_ram.memory[40][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11761_ (.D(_00283_),
    .CLK(net396),
    .Q(\u_cpu.rf_ram.memory[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11762_ (.D(_00284_),
    .CLK(net393),
    .Q(\u_cpu.rf_ram.memory[40][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11763_ (.D(_00285_),
    .CLK(net300),
    .Q(\u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11764_ (.D(_00286_),
    .CLK(net300),
    .Q(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11765_ (.D(_00287_),
    .CLK(net301),
    .Q(\u_cpu.rf_ram.memory[119][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00288_),
    .CLK(net345),
    .Q(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11767_ (.D(_00289_),
    .CLK(net345),
    .Q(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11768_ (.D(_00290_),
    .CLK(net394),
    .Q(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00291_),
    .CLK(net394),
    .Q(\u_cpu.rf_ram.memory[119][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00292_),
    .CLK(net393),
    .Q(\u_cpu.rf_ram.memory[119][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00293_),
    .CLK(net91),
    .Q(\u_cpu.rf_ram.memory[129][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00294_),
    .CLK(net91),
    .Q(\u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00295_),
    .CLK(net84),
    .Q(\u_cpu.rf_ram.memory[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00296_),
    .CLK(net91),
    .Q(\u_cpu.rf_ram.memory[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00297_),
    .CLK(net91),
    .Q(\u_cpu.rf_ram.memory[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00298_),
    .CLK(net84),
    .Q(\u_cpu.rf_ram.memory[129][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00299_),
    .CLK(net84),
    .Q(\u_cpu.rf_ram.memory[129][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00300_),
    .CLK(net85),
    .Q(\u_cpu.rf_ram.memory[129][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00301_),
    .CLK(net273),
    .Q(\u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00302_),
    .CLK(net268),
    .Q(\u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00303_),
    .CLK(net273),
    .Q(\u_cpu.rf_ram.memory[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00304_),
    .CLK(net269),
    .Q(\u_cpu.rf_ram.memory[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00305_),
    .CLK(net273),
    .Q(\u_cpu.rf_ram.memory[139][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00306_),
    .CLK(net274),
    .Q(\u_cpu.rf_ram.memory[139][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00307_),
    .CLK(net274),
    .Q(\u_cpu.rf_ram.memory[139][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00308_),
    .CLK(net268),
    .Q(\u_cpu.rf_ram.memory[139][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00309_),
    .CLK(net166),
    .Q(\u_cpu.rf_ram.memory[77][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00310_),
    .CLK(net166),
    .Q(\u_cpu.rf_ram.memory[77][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00311_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[77][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00312_),
    .CLK(net167),
    .Q(\u_cpu.rf_ram.memory[77][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00313_),
    .CLK(net167),
    .Q(\u_cpu.rf_ram.memory[77][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00314_),
    .CLK(net167),
    .Q(\u_cpu.rf_ram.memory[77][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00315_),
    .CLK(net167),
    .Q(\u_cpu.rf_ram.memory[77][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00316_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[77][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00317_),
    .CLK(net18),
    .Q(\u_cpu.rf_ram.memory[74][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00318_),
    .CLK(net34),
    .Q(\u_cpu.rf_ram.memory[74][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00319_),
    .CLK(net15),
    .Q(\u_cpu.rf_ram.memory[74][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00320_),
    .CLK(net15),
    .Q(\u_cpu.rf_ram.memory[74][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00321_),
    .CLK(net18),
    .Q(\u_cpu.rf_ram.memory[74][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00322_),
    .CLK(net34),
    .Q(\u_cpu.rf_ram.memory[74][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00323_),
    .CLK(net34),
    .Q(\u_cpu.rf_ram.memory[74][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00324_),
    .CLK(net34),
    .Q(\u_cpu.rf_ram.memory[74][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00325_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00326_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00327_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[76][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00328_),
    .CLK(net128),
    .Q(\u_cpu.rf_ram.memory[76][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00329_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[76][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00330_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[76][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00331_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[76][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00332_),
    .CLK(net126),
    .Q(\u_cpu.rf_ram.memory[76][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00333_),
    .CLK(net35),
    .Q(\u_cpu.rf_ram.memory[75][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11812_ (.D(_00334_),
    .CLK(net34),
    .Q(\u_cpu.rf_ram.memory[75][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11813_ (.D(_00335_),
    .CLK(net16),
    .Q(\u_cpu.rf_ram.memory[75][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11814_ (.D(_00336_),
    .CLK(net16),
    .Q(\u_cpu.rf_ram.memory[75][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00337_),
    .CLK(net18),
    .Q(\u_cpu.rf_ram.memory[75][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11816_ (.D(_00338_),
    .CLK(net35),
    .Q(\u_cpu.rf_ram.memory[75][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11817_ (.D(_00339_),
    .CLK(net35),
    .Q(\u_cpu.rf_ram.memory[75][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11818_ (.D(_00340_),
    .CLK(net35),
    .Q(\u_cpu.rf_ram.memory[75][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00341_),
    .CLK(net199),
    .Q(\u_cpu.rf_ram.memory[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11820_ (.D(_00342_),
    .CLK(net199),
    .Q(\u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11821_ (.D(_00343_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00344_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00345_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00346_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00347_),
    .CLK(net204),
    .Q(\u_cpu.rf_ram.memory[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00348_),
    .CLK(net199),
    .Q(\u_cpu.rf_ram.memory[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00349_),
    .CLK(net19),
    .Q(\u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00350_),
    .CLK(net18),
    .Q(\u_cpu.rf_ram.memory[68][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00351_),
    .CLK(net11),
    .Q(\u_cpu.rf_ram.memory[68][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11830_ (.D(_00352_),
    .CLK(net11),
    .Q(\u_cpu.rf_ram.memory[68][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00353_),
    .CLK(net11),
    .Q(\u_cpu.rf_ram.memory[68][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00354_),
    .CLK(net12),
    .Q(\u_cpu.rf_ram.memory[68][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00355_),
    .CLK(net12),
    .Q(\u_cpu.rf_ram.memory[68][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00356_),
    .CLK(net19),
    .Q(\u_cpu.rf_ram.memory[68][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00357_),
    .CLK(net105),
    .Q(\u_cpu.rf_ram.memory[67][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00358_),
    .CLK(net105),
    .Q(\u_cpu.rf_ram.memory[67][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00359_),
    .CLK(net97),
    .Q(\u_cpu.rf_ram.memory[67][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00360_),
    .CLK(net97),
    .Q(\u_cpu.rf_ram.memory[67][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00361_),
    .CLK(net97),
    .Q(\u_cpu.rf_ram.memory[67][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11840_ (.D(_00362_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[67][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11841_ (.D(_00363_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[67][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11842_ (.D(_00364_),
    .CLK(net106),
    .Q(\u_cpu.rf_ram.memory[67][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00365_),
    .CLK(net107),
    .Q(\u_cpu.rf_ram.memory[66][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00366_),
    .CLK(net107),
    .Q(\u_cpu.rf_ram.memory[66][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00367_),
    .CLK(net100),
    .Q(\u_cpu.rf_ram.memory[66][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00368_),
    .CLK(net100),
    .Q(\u_cpu.rf_ram.memory[66][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00369_),
    .CLK(net100),
    .Q(\u_cpu.rf_ram.memory[66][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11848_ (.D(_00370_),
    .CLK(net102),
    .Q(\u_cpu.rf_ram.memory[66][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11849_ (.D(_00371_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[66][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00372_),
    .CLK(net106),
    .Q(\u_cpu.rf_ram.memory[66][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00373_),
    .CLK(net105),
    .Q(\u_cpu.rf_ram.memory[65][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00374_),
    .CLK(net107),
    .Q(\u_cpu.rf_ram.memory[65][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00375_),
    .CLK(net97),
    .Q(\u_cpu.rf_ram.memory[65][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00376_),
    .CLK(net99),
    .Q(\u_cpu.rf_ram.memory[65][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00377_),
    .CLK(net97),
    .Q(\u_cpu.rf_ram.memory[65][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00378_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[65][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00379_),
    .CLK(net99),
    .Q(\u_cpu.rf_ram.memory[65][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00380_),
    .CLK(net106),
    .Q(\u_cpu.rf_ram.memory[65][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11859_ (.D(_00381_),
    .CLK(net108),
    .Q(\u_cpu.rf_ram.memory[64][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00382_),
    .CLK(net108),
    .Q(\u_cpu.rf_ram.memory[64][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00383_),
    .CLK(net102),
    .Q(\u_cpu.rf_ram.memory[64][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11862_ (.D(_00384_),
    .CLK(net102),
    .Q(\u_cpu.rf_ram.memory[64][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00385_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[64][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00386_),
    .CLK(net105),
    .Q(\u_cpu.rf_ram.memory[64][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00387_),
    .CLK(net105),
    .Q(\u_cpu.rf_ram.memory[64][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00388_),
    .CLK(net106),
    .Q(\u_cpu.rf_ram.memory[64][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00389_),
    .CLK(net183),
    .Q(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00390_),
    .CLK(net183),
    .Q(\u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00391_),
    .CLK(net166),
    .Q(\u_cpu.rf_ram.memory[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00392_),
    .CLK(net183),
    .Q(\u_cpu.rf_ram.memory[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00393_),
    .CLK(net168),
    .Q(\u_cpu.rf_ram.memory[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00394_),
    .CLK(net183),
    .Q(\u_cpu.rf_ram.memory[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11873_ (.D(_00395_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11874_ (.D(_00396_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11875_ (.D(_00397_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[63][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11876_ (.D(_00398_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[63][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11877_ (.D(_00399_),
    .CLK(net182),
    .Q(\u_cpu.rf_ram.memory[63][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00400_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00401_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00402_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[63][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00403_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[63][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00404_),
    .CLK(net167),
    .Q(\u_cpu.rf_ram.memory[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00405_),
    .CLK(net86),
    .Q(\u_cpu.rf_ram.memory[62][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00406_),
    .CLK(net86),
    .Q(\u_cpu.rf_ram.memory[62][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00407_),
    .CLK(net87),
    .Q(\u_cpu.rf_ram.memory[62][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00408_),
    .CLK(net89),
    .Q(\u_cpu.rf_ram.memory[62][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00409_),
    .CLK(net89),
    .Q(\u_cpu.rf_ram.memory[62][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00410_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11889_ (.D(_00411_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[62][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11890_ (.D(_00412_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[62][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11891_ (.D(_00413_),
    .CLK(net182),
    .Q(\u_cpu.rf_ram.memory[61][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11892_ (.D(_00414_),
    .CLK(net87),
    .Q(\u_cpu.rf_ram.memory[61][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11893_ (.D(_00415_),
    .CLK(net87),
    .Q(\u_cpu.rf_ram.memory[61][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11894_ (.D(_00416_),
    .CLK(net89),
    .Q(\u_cpu.rf_ram.memory[61][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11895_ (.D(_00417_),
    .CLK(net89),
    .Q(\u_cpu.rf_ram.memory[61][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11896_ (.D(_00418_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[61][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11897_ (.D(_00419_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[61][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11898_ (.D(_00420_),
    .CLK(net372),
    .Q(\u_cpu.rf_ram.memory[61][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11899_ (.D(_00421_),
    .CLK(net372),
    .Q(\u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00422_),
    .CLK(net89),
    .Q(\u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11901_ (.D(_00423_),
    .CLK(net90),
    .Q(\u_cpu.rf_ram.memory[60][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00424_),
    .CLK(net90),
    .Q(\u_cpu.rf_ram.memory[60][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00425_),
    .CLK(net90),
    .Q(\u_cpu.rf_ram.memory[60][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00426_),
    .CLK(net271),
    .Q(\u_cpu.rf_ram.memory[60][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00427_),
    .CLK(net271),
    .Q(\u_cpu.rf_ram.memory[60][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11906_ (.D(_00428_),
    .CLK(net271),
    .Q(\u_cpu.rf_ram.memory[60][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11907_ (.D(_00429_),
    .CLK(net375),
    .Q(\u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11908_ (.D(_00430_),
    .CLK(net275),
    .Q(\u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11909_ (.D(_00431_),
    .CLK(net275),
    .Q(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00432_),
    .CLK(net275),
    .Q(\u_cpu.rf_ram.memory[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00433_),
    .CLK(net276),
    .Q(\u_cpu.rf_ram.memory[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11912_ (.D(_00434_),
    .CLK(net276),
    .Q(\u_cpu.rf_ram.memory[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00435_),
    .CLK(net375),
    .Q(\u_cpu.rf_ram.memory[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00436_),
    .CLK(net375),
    .Q(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11915_ (.D(_00437_),
    .CLK(net213),
    .Q(\u_cpu.rf_ram.memory[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11916_ (.D(_00438_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11917_ (.D(_00439_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11918_ (.D(_00440_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11919_ (.D(_00441_),
    .CLK(net221),
    .Q(\u_cpu.rf_ram.memory[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00442_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00443_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00444_),
    .CLK(net213),
    .Q(\u_cpu.rf_ram.memory[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00445_),
    .CLK(net73),
    .Q(\u_cpu.rf_ram.memory[58][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11924_ (.D(_00446_),
    .CLK(net73),
    .Q(\u_cpu.rf_ram.memory[58][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11925_ (.D(_00447_),
    .CLK(net86),
    .Q(\u_cpu.rf_ram.memory[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11926_ (.D(_00448_),
    .CLK(net86),
    .Q(\u_cpu.rf_ram.memory[58][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11927_ (.D(_00449_),
    .CLK(net86),
    .Q(\u_cpu.rf_ram.memory[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11928_ (.D(_00450_),
    .CLK(net73),
    .Q(\u_cpu.rf_ram.memory[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11929_ (.D(_00451_),
    .CLK(net74),
    .Q(\u_cpu.rf_ram.memory[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11930_ (.D(_00452_),
    .CLK(net72),
    .Q(\u_cpu.rf_ram.memory[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00453_),
    .CLK(net70),
    .Q(\u_cpu.rf_ram.memory[57][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00454_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[57][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00455_),
    .CLK(net73),
    .Q(\u_cpu.rf_ram.memory[57][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00456_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram.memory[57][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00457_),
    .CLK(net69),
    .Q(\u_cpu.rf_ram.memory[57][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11936_ (.D(_00458_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[57][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11937_ (.D(_00459_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[57][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00460_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[57][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11939_ (.D(_00461_),
    .CLK(net68),
    .Q(\u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11940_ (.D(_00462_),
    .CLK(net68),
    .Q(\u_cpu.rf_ram.memory[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11941_ (.D(_00463_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram.memory[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11942_ (.D(_00464_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram.memory[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_00465_),
    .CLK(net69),
    .Q(\u_cpu.rf_ram.memory[56][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11944_ (.D(_00466_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11945_ (.D(_00467_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[56][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_00468_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[56][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_00469_),
    .CLK(net23),
    .Q(\u_cpu.rf_ram.memory[55][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11948_ (.D(_00470_),
    .CLK(net23),
    .Q(\u_cpu.rf_ram.memory[55][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11949_ (.D(_00471_),
    .CLK(net27),
    .Q(\u_cpu.rf_ram.memory[55][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11950_ (.D(_00472_),
    .CLK(net25),
    .Q(\u_cpu.rf_ram.memory[55][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11951_ (.D(_00473_),
    .CLK(net25),
    .Q(\u_cpu.rf_ram.memory[55][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_00474_),
    .CLK(net25),
    .Q(\u_cpu.rf_ram.memory[55][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_00475_),
    .CLK(net25),
    .Q(\u_cpu.rf_ram.memory[55][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11954_ (.D(_00476_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[55][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_00477_),
    .CLK(net23),
    .Q(\u_cpu.rf_ram.memory[54][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11956_ (.D(_00478_),
    .CLK(net23),
    .Q(\u_cpu.rf_ram.memory[54][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11957_ (.D(_00479_),
    .CLK(net23),
    .Q(\u_cpu.rf_ram.memory[54][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_00480_),
    .CLK(net24),
    .Q(\u_cpu.rf_ram.memory[54][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_00481_),
    .CLK(net24),
    .Q(\u_cpu.rf_ram.memory[54][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11960_ (.D(_00482_),
    .CLK(net24),
    .Q(\u_cpu.rf_ram.memory[54][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11961_ (.D(_00483_),
    .CLK(net24),
    .Q(\u_cpu.rf_ram.memory[54][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11962_ (.D(_00484_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[54][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11963_ (.D(_00485_),
    .CLK(net28),
    .Q(\u_cpu.rf_ram.memory[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11964_ (.D(_00486_),
    .CLK(net28),
    .Q(\u_cpu.rf_ram.memory[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_00487_),
    .CLK(net28),
    .Q(\u_cpu.rf_ram.memory[53][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_00488_),
    .CLK(net30),
    .Q(\u_cpu.rf_ram.memory[53][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_00489_),
    .CLK(net30),
    .Q(\u_cpu.rf_ram.memory[53][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_00490_),
    .CLK(net30),
    .Q(\u_cpu.rf_ram.memory[53][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11969_ (.D(_00491_),
    .CLK(net31),
    .Q(\u_cpu.rf_ram.memory[53][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_00492_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[53][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11971_ (.D(_00493_),
    .CLK(net28),
    .Q(\u_cpu.rf_ram.memory[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11972_ (.D(_00494_),
    .CLK(net28),
    .Q(\u_cpu.rf_ram.memory[52][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11973_ (.D(_00495_),
    .CLK(net29),
    .Q(\u_cpu.rf_ram.memory[52][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11974_ (.D(_00496_),
    .CLK(net29),
    .Q(\u_cpu.rf_ram.memory[52][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11975_ (.D(_00497_),
    .CLK(net31),
    .Q(\u_cpu.rf_ram.memory[52][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11976_ (.D(_00498_),
    .CLK(net58),
    .Q(\u_cpu.rf_ram.memory[52][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11977_ (.D(_00499_),
    .CLK(net58),
    .Q(\u_cpu.rf_ram.memory[52][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11978_ (.D(_00500_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[52][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11979_ (.D(_00501_),
    .CLK(net221),
    .Q(\u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11980_ (.D(_00502_),
    .CLK(net221),
    .Q(\u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11981_ (.D(_00503_),
    .CLK(net421),
    .Q(\u_cpu.rf_ram.memory[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11982_ (.D(_00504_),
    .CLK(net421),
    .Q(\u_cpu.rf_ram.memory[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11983_ (.D(_00505_),
    .CLK(net421),
    .Q(\u_cpu.rf_ram.memory[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11984_ (.D(_00506_),
    .CLK(net221),
    .Q(\u_cpu.rf_ram.memory[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11985_ (.D(_00507_),
    .CLK(net214),
    .Q(\u_cpu.rf_ram.memory[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11986_ (.D(_00508_),
    .CLK(net214),
    .Q(\u_cpu.rf_ram.memory[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11987_ (.D(_00509_),
    .CLK(net223),
    .Q(\u_cpu.rf_ram.memory[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11988_ (.D(_00510_),
    .CLK(net223),
    .Q(\u_cpu.rf_ram.memory[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11989_ (.D(_00511_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11990_ (.D(_00512_),
    .CLK(net420),
    .Q(\u_cpu.rf_ram.memory[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11991_ (.D(_00513_),
    .CLK(net420),
    .Q(\u_cpu.rf_ram.memory[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11992_ (.D(_00514_),
    .CLK(net223),
    .Q(\u_cpu.rf_ram.memory[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11993_ (.D(_00515_),
    .CLK(net223),
    .Q(\u_cpu.rf_ram.memory[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11994_ (.D(_00516_),
    .CLK(net223),
    .Q(\u_cpu.rf_ram.memory[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_00000_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11996_ (.D(_00001_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_00002_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_00003_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11999_ (.D(_00004_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_00005_),
    .CLK(net292),
    .Q(\u_cpu.rf_ram.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_00006_),
    .CLK(net292),
    .Q(\u_cpu.rf_ram.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_00007_),
    .CLK(net283),
    .Q(\u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12003_ (.D(_00517_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[142][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12004_ (.D(_00518_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[142][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12005_ (.D(_00519_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[142][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12006_ (.D(_00520_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[142][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12007_ (.D(_00521_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[142][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12008_ (.D(_00522_),
    .CLK(net58),
    .Q(\u_cpu.rf_ram.memory[142][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(_00523_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[142][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12010_ (.D(_00524_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[142][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(_00525_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[141][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(_00526_),
    .CLK(net61),
    .Q(\u_cpu.rf_ram.memory[141][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(_00527_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[141][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12014_ (.D(_00528_),
    .CLK(net43),
    .Q(\u_cpu.rf_ram.memory[141][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12015_ (.D(_00529_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[141][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12016_ (.D(_00530_),
    .CLK(net57),
    .Q(\u_cpu.rf_ram.memory[141][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12017_ (.D(_00531_),
    .CLK(net61),
    .Q(\u_cpu.rf_ram.memory[141][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12018_ (.D(_00532_),
    .CLK(net69),
    .Q(\u_cpu.rf_ram.memory[141][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12019_ (.D(_00533_),
    .CLK(net57),
    .Q(\u_cpu.rf_ram.memory[140][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12020_ (.D(_00534_),
    .CLK(net61),
    .Q(\u_cpu.rf_ram.memory[140][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12021_ (.D(_00535_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[140][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12022_ (.D(_00536_),
    .CLK(net43),
    .Q(\u_cpu.rf_ram.memory[140][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12023_ (.D(_00537_),
    .CLK(net43),
    .Q(\u_cpu.rf_ram.memory[140][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12024_ (.D(_00538_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[140][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12025_ (.D(_00539_),
    .CLK(net61),
    .Q(\u_cpu.rf_ram.memory[140][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12026_ (.D(_00540_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram.memory[140][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12027_ (.D(_00541_),
    .CLK(net224),
    .Q(\u_cpu.rf_ram.memory[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12028_ (.D(_00542_),
    .CLK(net224),
    .Q(\u_cpu.rf_ram.memory[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12029_ (.D(_00543_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12030_ (.D(_00544_),
    .CLK(net420),
    .Q(\u_cpu.rf_ram.memory[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12031_ (.D(_00545_),
    .CLK(net420),
    .Q(\u_cpu.rf_ram.memory[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12032_ (.D(_00546_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12033_ (.D(_00547_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12034_ (.D(_00548_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12035_ (.D(_00549_),
    .CLK(net24),
    .Q(\u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12036_ (.D(_00550_),
    .CLK(net26),
    .Q(\u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(_00551_),
    .CLK(net22),
    .Q(\u_cpu.rf_ram.memory[72][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12038_ (.D(_00552_),
    .CLK(net22),
    .Q(\u_cpu.rf_ram.memory[72][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12039_ (.D(_00553_),
    .CLK(net22),
    .Q(\u_cpu.rf_ram.memory[72][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12040_ (.D(_00554_),
    .CLK(net25),
    .Q(\u_cpu.rf_ram.memory[72][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12041_ (.D(_00555_),
    .CLK(net26),
    .Q(\u_cpu.rf_ram.memory[72][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(_00556_),
    .CLK(net33),
    .Q(\u_cpu.rf_ram.memory[72][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12043_ (.D(_00557_),
    .CLK(net33),
    .Q(\u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12044_ (.D(_00558_),
    .CLK(net33),
    .Q(\u_cpu.rf_ram.memory[73][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12045_ (.D(_00559_),
    .CLK(net16),
    .Q(\u_cpu.rf_ram.memory[73][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12046_ (.D(_00560_),
    .CLK(net17),
    .Q(\u_cpu.rf_ram.memory[73][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12047_ (.D(_00561_),
    .CLK(net17),
    .Q(\u_cpu.rf_ram.memory[73][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12048_ (.D(_00562_),
    .CLK(net33),
    .Q(\u_cpu.rf_ram.memory[73][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12049_ (.D(_00563_),
    .CLK(net33),
    .Q(\u_cpu.rf_ram.memory[73][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(_00564_),
    .CLK(net36),
    .Q(\u_cpu.rf_ram.memory[73][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12051_ (.D(_00565_),
    .CLK(net15),
    .Q(\u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12052_ (.D(_00566_),
    .CLK(net9),
    .Q(\u_cpu.rf_ram.memory[71][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12053_ (.D(_00567_),
    .CLK(net8),
    .Q(\u_cpu.rf_ram.memory[71][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12054_ (.D(_00568_),
    .CLK(net8),
    .Q(\u_cpu.rf_ram.memory[71][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12055_ (.D(_00569_),
    .CLK(net9),
    .Q(\u_cpu.rf_ram.memory[71][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12056_ (.D(_00570_),
    .CLK(net9),
    .Q(\u_cpu.rf_ram.memory[71][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12057_ (.D(_00571_),
    .CLK(net9),
    .Q(\u_cpu.rf_ram.memory[71][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12058_ (.D(_00572_),
    .CLK(net16),
    .Q(\u_cpu.rf_ram.memory[71][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12059_ (.D(_00573_),
    .CLK(net15),
    .Q(\u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12060_ (.D(_00574_),
    .CLK(net22),
    .Q(\u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12061_ (.D(_00575_),
    .CLK(net8),
    .Q(\u_cpu.rf_ram.memory[70][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12062_ (.D(_00576_),
    .CLK(net8),
    .Q(\u_cpu.rf_ram.memory[70][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12063_ (.D(_00577_),
    .CLK(net8),
    .Q(\u_cpu.rf_ram.memory[70][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12064_ (.D(_00578_),
    .CLK(net10),
    .Q(\u_cpu.rf_ram.memory[70][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12065_ (.D(_00579_),
    .CLK(net10),
    .Q(\u_cpu.rf_ram.memory[70][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12066_ (.D(_00580_),
    .CLK(net15),
    .Q(\u_cpu.rf_ram.memory[70][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12067_ (.D(_00581_),
    .CLK(net58),
    .Q(\u_cpu.rf_ram.memory[143][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12068_ (.D(_00582_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[143][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12069_ (.D(_00583_),
    .CLK(net58),
    .Q(\u_cpu.rf_ram.memory[143][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12070_ (.D(_00584_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[143][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12071_ (.D(_00585_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[143][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12072_ (.D(_00586_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[143][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12073_ (.D(_00587_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[143][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12074_ (.D(_00588_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[143][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12075_ (.D(_00589_),
    .CLK(net222),
    .Q(\u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12076_ (.D(_00590_),
    .CLK(net219),
    .Q(\u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12077_ (.D(_00591_),
    .CLK(net222),
    .Q(\u_cpu.rf_ram.memory[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12078_ (.D(_00592_),
    .CLK(net225),
    .Q(\u_cpu.rf_ram.memory[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12079_ (.D(_00593_),
    .CLK(net227),
    .Q(\u_cpu.rf_ram.memory[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12080_ (.D(_00594_),
    .CLK(net222),
    .Q(\u_cpu.rf_ram.memory[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12081_ (.D(_00595_),
    .CLK(net222),
    .Q(\u_cpu.rf_ram.memory[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12082_ (.D(_00596_),
    .CLK(net222),
    .Q(\u_cpu.rf_ram.memory[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12083_ (.D(_00597_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12084_ (.D(_00598_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12085_ (.D(_00599_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12086_ (.D(_00600_),
    .CLK(net64),
    .Q(\u_cpu.rf_ram.memory[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12087_ (.D(_00601_),
    .CLK(net64),
    .Q(\u_cpu.rf_ram.memory[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12088_ (.D(_00602_),
    .CLK(net72),
    .Q(\u_cpu.rf_ram.memory[138][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12089_ (.D(_00603_),
    .CLK(net72),
    .Q(\u_cpu.rf_ram.memory[138][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12090_ (.D(_00604_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram.memory[138][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12091_ (.D(_00605_),
    .CLK(net337),
    .Q(\u_cpu.rf_ram.memory[39][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12092_ (.D(_00606_),
    .CLK(net337),
    .Q(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12093_ (.D(_00607_),
    .CLK(net336),
    .Q(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12094_ (.D(_00608_),
    .CLK(net337),
    .Q(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12095_ (.D(_00609_),
    .CLK(net336),
    .Q(\u_cpu.rf_ram.memory[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12096_ (.D(_00610_),
    .CLK(net338),
    .Q(\u_cpu.rf_ram.memory[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12097_ (.D(_00611_),
    .CLK(net343),
    .Q(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12098_ (.D(_00612_),
    .CLK(net344),
    .Q(\u_cpu.rf_ram.memory[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12099_ (.D(_00613_),
    .CLK(net264),
    .Q(\u_cpu.rf_ram.memory[137][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12100_ (.D(_00614_),
    .CLK(net260),
    .Q(\u_cpu.rf_ram.memory[137][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12101_ (.D(_00615_),
    .CLK(net264),
    .Q(\u_cpu.rf_ram.memory[137][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12102_ (.D(_00616_),
    .CLK(net261),
    .Q(\u_cpu.rf_ram.memory[137][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12103_ (.D(_00617_),
    .CLK(net264),
    .Q(\u_cpu.rf_ram.memory[137][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12104_ (.D(_00618_),
    .CLK(net273),
    .Q(\u_cpu.rf_ram.memory[137][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12105_ (.D(_00619_),
    .CLK(net269),
    .Q(\u_cpu.rf_ram.memory[137][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12106_ (.D(_00620_),
    .CLK(net273),
    .Q(\u_cpu.rf_ram.memory[137][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12107_ (.D(_00621_),
    .CLK(net281),
    .Q(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12108_ (.D(_00622_),
    .CLK(net282),
    .Q(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12109_ (.D(_00623_),
    .CLK(net293),
    .Q(\u_cpu.rf_ram.memory[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12110_ (.D(_00624_),
    .CLK(net293),
    .Q(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12111_ (.D(_00625_),
    .CLK(net282),
    .Q(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12112_ (.D(_00626_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12113_ (.D(_00627_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12114_ (.D(_00628_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.memory[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12115_ (.D(_00629_),
    .CLK(net264),
    .Q(\u_cpu.rf_ram.memory[136][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12116_ (.D(_00630_),
    .CLK(net264),
    .Q(\u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12117_ (.D(_00631_),
    .CLK(net265),
    .Q(\u_cpu.rf_ram.memory[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12118_ (.D(_00632_),
    .CLK(net265),
    .Q(\u_cpu.rf_ram.memory[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12119_ (.D(_00633_),
    .CLK(net283),
    .Q(\u_cpu.rf_ram.memory[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12120_ (.D(_00634_),
    .CLK(net274),
    .Q(\u_cpu.rf_ram.memory[136][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12121_ (.D(_00635_),
    .CLK(net274),
    .Q(\u_cpu.rf_ram.memory[136][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12122_ (.D(_00636_),
    .CLK(net265),
    .Q(\u_cpu.rf_ram.memory[136][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12123_ (.D(_00637_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[135][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12124_ (.D(_00638_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[135][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12125_ (.D(_00639_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[135][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12126_ (.D(_00640_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[135][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12127_ (.D(_00641_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[135][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12128_ (.D(_00642_),
    .CLK(net259),
    .Q(\u_cpu.rf_ram.memory[135][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12129_ (.D(_00643_),
    .CLK(net259),
    .Q(\u_cpu.rf_ram.memory[135][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12130_ (.D(_00644_),
    .CLK(net259),
    .Q(\u_cpu.rf_ram.memory[135][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12131_ (.D(_00645_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[134][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12132_ (.D(_00646_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[134][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12133_ (.D(_00647_),
    .CLK(net61),
    .Q(\u_cpu.rf_ram.memory[134][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12134_ (.D(_00648_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[134][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12135_ (.D(_00649_),
    .CLK(net43),
    .Q(\u_cpu.rf_ram.memory[134][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12136_ (.D(_00650_),
    .CLK(net62),
    .Q(\u_cpu.rf_ram.memory[134][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12137_ (.D(_00651_),
    .CLK(net62),
    .Q(\u_cpu.rf_ram.memory[134][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12138_ (.D(_00652_),
    .CLK(net82),
    .Q(\u_cpu.rf_ram.memory[134][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12139_ (.D(_00653_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[133][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12140_ (.D(_00654_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram.memory[133][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12141_ (.D(_00655_),
    .CLK(net43),
    .Q(\u_cpu.rf_ram.memory[133][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12142_ (.D(_00656_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[133][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12143_ (.D(_00657_),
    .CLK(net44),
    .Q(\u_cpu.rf_ram.memory[133][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12144_ (.D(_00658_),
    .CLK(net62),
    .Q(\u_cpu.rf_ram.memory[133][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12145_ (.D(_00659_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[133][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12146_ (.D(_00660_),
    .CLK(net82),
    .Q(\u_cpu.rf_ram.memory[133][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12147_ (.D(_00661_),
    .CLK(net78),
    .Q(\u_cpu.rf_ram.memory[132][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12148_ (.D(_00662_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram.memory[132][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12149_ (.D(_00663_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[132][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12150_ (.D(_00664_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram.memory[132][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12151_ (.D(_00665_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[132][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12152_ (.D(_00666_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[132][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12153_ (.D(_00667_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[132][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12154_ (.D(_00668_),
    .CLK(net82),
    .Q(\u_cpu.rf_ram.memory[132][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12155_ (.D(_00669_),
    .CLK(net80),
    .Q(\u_cpu.rf_ram.memory[131][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12156_ (.D(_00670_),
    .CLK(net82),
    .Q(\u_cpu.rf_ram.memory[131][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12157_ (.D(_00671_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[131][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12158_ (.D(_00672_),
    .CLK(net78),
    .Q(\u_cpu.rf_ram.memory[131][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12159_ (.D(_00673_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[131][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12160_ (.D(_00674_),
    .CLK(net84),
    .Q(\u_cpu.rf_ram.memory[131][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12161_ (.D(_00675_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[131][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12162_ (.D(_00676_),
    .CLK(net85),
    .Q(\u_cpu.rf_ram.memory[131][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12163_ (.D(_00677_),
    .CLK(net82),
    .Q(\u_cpu.rf_ram.memory[130][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12164_ (.D(_00678_),
    .CLK(net83),
    .Q(\u_cpu.rf_ram.memory[130][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12165_ (.D(_00679_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[130][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12166_ (.D(_00680_),
    .CLK(net80),
    .Q(\u_cpu.rf_ram.memory[130][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12167_ (.D(_00681_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[130][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12168_ (.D(_00682_),
    .CLK(net84),
    .Q(\u_cpu.rf_ram.memory[130][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12169_ (.D(_00683_),
    .CLK(net80),
    .Q(\u_cpu.rf_ram.memory[130][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12170_ (.D(_00684_),
    .CLK(net85),
    .Q(\u_cpu.rf_ram.memory[130][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12171_ (.D(_00685_),
    .CLK(net424),
    .Q(\u_cpu.rf_ram.memory[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12172_ (.D(_00686_),
    .CLK(net425),
    .Q(\u_cpu.rf_ram.memory[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12173_ (.D(_00687_),
    .CLK(net424),
    .Q(\u_cpu.rf_ram.memory[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12174_ (.D(_00688_),
    .CLK(net424),
    .Q(\u_cpu.rf_ram.memory[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12175_ (.D(_00689_),
    .CLK(net424),
    .Q(\u_cpu.rf_ram.memory[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12176_ (.D(_00690_),
    .CLK(net425),
    .Q(\u_cpu.rf_ram.memory[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12177_ (.D(_00691_),
    .CLK(net425),
    .Q(\u_cpu.rf_ram.memory[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12178_ (.D(_00692_),
    .CLK(net424),
    .Q(\u_cpu.rf_ram.memory[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12179_ (.D(_00693_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12180_ (.D(_00694_),
    .CLK(net192),
    .Q(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12181_ (.D(_00695_),
    .CLK(net374),
    .Q(\u_cpu.rf_ram.memory[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12182_ (.D(_00696_),
    .CLK(net372),
    .Q(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12183_ (.D(_00697_),
    .CLK(net373),
    .Q(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12184_ (.D(_00698_),
    .CLK(net372),
    .Q(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12185_ (.D(_00699_),
    .CLK(net372),
    .Q(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12186_ (.D(_00700_),
    .CLK(net373),
    .Q(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12187_ (.D(_00701_),
    .CLK(net260),
    .Q(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12188_ (.D(_00702_),
    .CLK(net260),
    .Q(\u_cpu.rf_ram.memory[128][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12189_ (.D(_00703_),
    .CLK(net261),
    .Q(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12190_ (.D(_00704_),
    .CLK(net260),
    .Q(\u_cpu.rf_ram.memory[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12191_ (.D(_00705_),
    .CLK(net260),
    .Q(\u_cpu.rf_ram.memory[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12192_ (.D(_00706_),
    .CLK(net268),
    .Q(\u_cpu.rf_ram.memory[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12193_ (.D(_00707_),
    .CLK(net268),
    .Q(\u_cpu.rf_ram.memory[128][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12194_ (.D(_00708_),
    .CLK(net268),
    .Q(\u_cpu.rf_ram.memory[128][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12195_ (.D(_00709_),
    .CLK(net293),
    .Q(\u_cpu.rf_ram.memory[127][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12196_ (.D(_00710_),
    .CLK(net296),
    .Q(\u_cpu.rf_ram.memory[127][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12197_ (.D(_00711_),
    .CLK(net298),
    .Q(\u_cpu.rf_ram.memory[127][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12198_ (.D(_00712_),
    .CLK(net298),
    .Q(\u_cpu.rf_ram.memory[127][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12199_ (.D(_00713_),
    .CLK(net343),
    .Q(\u_cpu.rf_ram.memory[127][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12200_ (.D(_00714_),
    .CLK(net345),
    .Q(\u_cpu.rf_ram.memory[127][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12201_ (.D(_00715_),
    .CLK(net345),
    .Q(\u_cpu.rf_ram.memory[127][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12202_ (.D(_00716_),
    .CLK(net300),
    .Q(\u_cpu.rf_ram.memory[127][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12203_ (.D(_00717_),
    .CLK(net296),
    .Q(\u_cpu.rf_ram.memory[126][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12204_ (.D(_00718_),
    .CLK(net296),
    .Q(\u_cpu.rf_ram.memory[126][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12205_ (.D(_00719_),
    .CLK(net298),
    .Q(\u_cpu.rf_ram.memory[126][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12206_ (.D(_00720_),
    .CLK(net298),
    .Q(\u_cpu.rf_ram.memory[126][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12207_ (.D(_00721_),
    .CLK(net299),
    .Q(\u_cpu.rf_ram.memory[126][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12208_ (.D(_00722_),
    .CLK(net301),
    .Q(\u_cpu.rf_ram.memory[126][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12209_ (.D(_00723_),
    .CLK(net301),
    .Q(\u_cpu.rf_ram.memory[126][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12210_ (.D(_00724_),
    .CLK(net300),
    .Q(\u_cpu.rf_ram.memory[126][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12211_ (.D(_00725_),
    .CLK(net294),
    .Q(\u_cpu.rf_ram.memory[125][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12212_ (.D(_00726_),
    .CLK(net294),
    .Q(\u_cpu.rf_ram.memory[125][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12213_ (.D(_00727_),
    .CLK(net298),
    .Q(\u_cpu.rf_ram.memory[125][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12214_ (.D(_00728_),
    .CLK(net299),
    .Q(\u_cpu.rf_ram.memory[125][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12215_ (.D(_00729_),
    .CLK(net343),
    .Q(\u_cpu.rf_ram.memory[125][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12216_ (.D(_00730_),
    .CLK(net343),
    .Q(\u_cpu.rf_ram.memory[125][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12217_ (.D(_00731_),
    .CLK(net343),
    .Q(\u_cpu.rf_ram.memory[125][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12218_ (.D(_00732_),
    .CLK(net300),
    .Q(\u_cpu.rf_ram.memory[125][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12219_ (.D(_00733_),
    .CLK(net348),
    .Q(\u_cpu.rf_ram.memory[124][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12220_ (.D(_00734_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[124][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12221_ (.D(_00735_),
    .CLK(net348),
    .Q(\u_cpu.rf_ram.memory[124][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12222_ (.D(_00736_),
    .CLK(net344),
    .Q(\u_cpu.rf_ram.memory[124][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12223_ (.D(_00737_),
    .CLK(net344),
    .Q(\u_cpu.rf_ram.memory[124][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12224_ (.D(_00738_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[124][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12225_ (.D(_00739_),
    .CLK(net345),
    .Q(\u_cpu.rf_ram.memory[124][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12226_ (.D(_00740_),
    .CLK(net346),
    .Q(\u_cpu.rf_ram.memory[124][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12227_ (.D(_00015_),
    .CLK(net287),
    .Q(\u_cpu.rf_ram_if.rdata1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12228_ (.D(_00016_),
    .CLK(net287),
    .Q(\u_cpu.rf_ram_if.rdata1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12229_ (.D(_00017_),
    .CLK(net287),
    .Q(\u_cpu.rf_ram_if.rdata1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12230_ (.D(_00018_),
    .CLK(net287),
    .Q(\u_cpu.rf_ram_if.rdata1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12231_ (.D(_00019_),
    .CLK(net281),
    .Q(\u_cpu.rf_ram_if.rdata1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12232_ (.D(_00020_),
    .CLK(net281),
    .Q(\u_cpu.rf_ram_if.rdata1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12233_ (.D(_00008_),
    .CLK(net285),
    .Q(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12234_ (.D(_00009_),
    .CLK(net285),
    .Q(\u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12235_ (.D(_00010_),
    .CLK(net287),
    .Q(\u_cpu.rf_ram_if.rdata0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12236_ (.D(_00011_),
    .CLK(net280),
    .Q(\u_cpu.rf_ram_if.rdata0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12237_ (.D(_00012_),
    .CLK(net279),
    .Q(\u_cpu.rf_ram_if.rdata0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12238_ (.D(_00013_),
    .CLK(net281),
    .Q(\u_cpu.rf_ram_if.rdata0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12239_ (.D(_00014_),
    .CLK(net279),
    .Q(\u_cpu.rf_ram_if.rdata0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12240_ (.D(_00741_),
    .CLK(net361),
    .Q(\u_cpu.rf_ram.memory[123][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12241_ (.D(_00742_),
    .CLK(net361),
    .Q(\u_cpu.rf_ram.memory[123][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12242_ (.D(_00743_),
    .CLK(net358),
    .Q(\u_cpu.rf_ram.memory[123][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12243_ (.D(_00744_),
    .CLK(net358),
    .Q(\u_cpu.rf_ram.memory[123][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12244_ (.D(_00745_),
    .CLK(net358),
    .Q(\u_cpu.rf_ram.memory[123][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12245_ (.D(_00746_),
    .CLK(net362),
    .Q(\u_cpu.rf_ram.memory[123][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12246_ (.D(_00747_),
    .CLK(net362),
    .Q(\u_cpu.rf_ram.memory[123][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12247_ (.D(_00748_),
    .CLK(net361),
    .Q(\u_cpu.rf_ram.memory[123][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12248_ (.D(_00749_),
    .CLK(net348),
    .Q(\u_cpu.rf_ram.memory[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12249_ (.D(_00750_),
    .CLK(net348),
    .Q(\u_cpu.rf_ram.memory[38][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12250_ (.D(_00751_),
    .CLK(net339),
    .Q(\u_cpu.rf_ram.memory[38][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12251_ (.D(_00752_),
    .CLK(net339),
    .Q(\u_cpu.rf_ram.memory[38][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12252_ (.D(_00753_),
    .CLK(net339),
    .Q(\u_cpu.rf_ram.memory[38][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12253_ (.D(_00754_),
    .CLK(net348),
    .Q(\u_cpu.rf_ram.memory[38][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12254_ (.D(_00755_),
    .CLK(net349),
    .Q(\u_cpu.rf_ram.memory[38][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12255_ (.D(_00756_),
    .CLK(net349),
    .Q(\u_cpu.rf_ram.memory[38][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12256_ (.D(_00757_),
    .CLK(net349),
    .Q(\u_cpu.rf_ram.memory[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12257_ (.D(_00758_),
    .CLK(net360),
    .Q(\u_cpu.rf_ram.memory[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12258_ (.D(_00759_),
    .CLK(net355),
    .Q(\u_cpu.rf_ram.memory[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12259_ (.D(_00760_),
    .CLK(net355),
    .Q(\u_cpu.rf_ram.memory[37][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12260_ (.D(_00761_),
    .CLK(net355),
    .Q(\u_cpu.rf_ram.memory[37][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12261_ (.D(_00762_),
    .CLK(net360),
    .Q(\u_cpu.rf_ram.memory[37][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12262_ (.D(_00763_),
    .CLK(net360),
    .Q(\u_cpu.rf_ram.memory[37][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12263_ (.D(_00764_),
    .CLK(net360),
    .Q(\u_cpu.rf_ram.memory[37][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12264_ (.D(_00765_),
    .CLK(net355),
    .Q(\u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12265_ (.D(_00766_),
    .CLK(net358),
    .Q(\u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12266_ (.D(_00767_),
    .CLK(net355),
    .Q(\u_cpu.rf_ram.memory[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12267_ (.D(_00768_),
    .CLK(net356),
    .Q(\u_cpu.rf_ram.memory[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12268_ (.D(_00769_),
    .CLK(net356),
    .Q(\u_cpu.rf_ram.memory[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12269_ (.D(_00770_),
    .CLK(net358),
    .Q(\u_cpu.rf_ram.memory[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12270_ (.D(_00771_),
    .CLK(net359),
    .Q(\u_cpu.rf_ram.memory[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12271_ (.D(_00772_),
    .CLK(net359),
    .Q(\u_cpu.rf_ram.memory[36][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12272_ (.D(_00773_),
    .CLK(net255),
    .Q(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12273_ (.D(_00774_),
    .CLK(net316),
    .Q(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12274_ (.D(_00775_),
    .CLK(net314),
    .Q(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12275_ (.D(_00776_),
    .CLK(net314),
    .Q(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12276_ (.D(_00777_),
    .CLK(net316),
    .Q(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12277_ (.D(_00778_),
    .CLK(net319),
    .Q(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12278_ (.D(_00779_),
    .CLK(net313),
    .Q(\u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12279_ (.D(_00780_),
    .CLK(net313),
    .Q(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12280_ (.D(_00781_),
    .CLK(net380),
    .Q(\u_cpu.rf_ram.memory[91][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12281_ (.D(_00782_),
    .CLK(net380),
    .Q(\u_cpu.rf_ram.memory[91][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12282_ (.D(_00783_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[91][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12283_ (.D(_00784_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[91][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12284_ (.D(_00785_),
    .CLK(net399),
    .Q(\u_cpu.rf_ram.memory[91][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12285_ (.D(_00786_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[91][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12286_ (.D(_00787_),
    .CLK(net399),
    .Q(\u_cpu.rf_ram.memory[91][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12287_ (.D(_00788_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[91][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12288_ (.D(_00789_),
    .CLK(net380),
    .Q(\u_cpu.rf_ram.memory[90][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12289_ (.D(_00790_),
    .CLK(net380),
    .Q(\u_cpu.rf_ram.memory[90][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12290_ (.D(_00791_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[90][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12291_ (.D(_00792_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[90][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12292_ (.D(_00793_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[90][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12293_ (.D(_00794_),
    .CLK(net380),
    .Q(\u_cpu.rf_ram.memory[90][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12294_ (.D(_00795_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[90][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12295_ (.D(_00796_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[90][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12296_ (.D(_00797_),
    .CLK(net314),
    .Q(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12297_ (.D(_00798_),
    .CLK(net255),
    .Q(\u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12298_ (.D(_00799_),
    .CLK(net315),
    .Q(\u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12299_ (.D(_00800_),
    .CLK(net316),
    .Q(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12300_ (.D(_00801_),
    .CLK(net315),
    .Q(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12301_ (.D(_00802_),
    .CLK(net197),
    .Q(\u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12302_ (.D(_00803_),
    .CLK(net207),
    .Q(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12303_ (.D(_00804_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12304_ (.D(_00805_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[92][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12305_ (.D(_00806_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[92][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12306_ (.D(_00807_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[92][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12307_ (.D(_00808_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[92][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12308_ (.D(_00809_),
    .CLK(net197),
    .Q(\u_cpu.rf_ram.memory[92][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12309_ (.D(_00810_),
    .CLK(net487),
    .Q(\u_cpu.rf_ram.memory[35][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12310_ (.D(_00811_),
    .CLK(net467),
    .Q(\u_cpu.rf_ram.memory[35][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12311_ (.D(_00812_),
    .CLK(net487),
    .Q(\u_cpu.rf_ram.memory[35][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12312_ (.D(_00813_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[35][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12313_ (.D(_00814_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[35][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12314_ (.D(_00815_),
    .CLK(net464),
    .Q(\u_cpu.rf_ram.memory[35][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12315_ (.D(_00816_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[35][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12316_ (.D(_00817_),
    .CLK(net465),
    .Q(\u_cpu.rf_ram.memory[35][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12317_ (.D(_00818_),
    .CLK(net487),
    .Q(\u_cpu.rf_ram.memory[34][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12318_ (.D(_00819_),
    .CLK(net467),
    .Q(\u_cpu.rf_ram.memory[34][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12319_ (.D(_00820_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[34][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12320_ (.D(_00821_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[34][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12321_ (.D(_00822_),
    .CLK(net487),
    .Q(\u_cpu.rf_ram.memory[34][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12322_ (.D(_00823_),
    .CLK(net467),
    .Q(\u_cpu.rf_ram.memory[34][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12323_ (.D(_00824_),
    .CLK(net487),
    .Q(\u_cpu.rf_ram.memory[34][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12324_ (.D(_00825_),
    .CLK(net468),
    .Q(\u_cpu.rf_ram.memory[34][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12325_ (.D(_00826_),
    .CLK(net454),
    .Q(\u_cpu.rf_ram.memory[117][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12326_ (.D(_00827_),
    .CLK(net351),
    .Q(\u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12327_ (.D(_00828_),
    .CLK(net361),
    .Q(\u_cpu.rf_ram.memory[117][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12328_ (.D(_00829_),
    .CLK(net351),
    .Q(\u_cpu.rf_ram.memory[117][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12329_ (.D(_00830_),
    .CLK(net351),
    .Q(\u_cpu.rf_ram.memory[117][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12330_ (.D(_00831_),
    .CLK(net454),
    .Q(\u_cpu.rf_ram.memory[117][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12331_ (.D(_00832_),
    .CLK(net454),
    .Q(\u_cpu.rf_ram.memory[117][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12332_ (.D(_00833_),
    .CLK(net454),
    .Q(\u_cpu.rf_ram.memory[117][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12333_ (.D(_00834_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[120][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12334_ (.D(_00835_),
    .CLK(net364),
    .Q(\u_cpu.rf_ram.memory[120][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12335_ (.D(_00836_),
    .CLK(net364),
    .Q(\u_cpu.rf_ram.memory[120][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12336_ (.D(_00837_),
    .CLK(net365),
    .Q(\u_cpu.rf_ram.memory[120][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12337_ (.D(_00838_),
    .CLK(net365),
    .Q(\u_cpu.rf_ram.memory[120][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12338_ (.D(_00839_),
    .CLK(net365),
    .Q(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12339_ (.D(_00840_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[120][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12340_ (.D(_00841_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[120][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12341_ (.D(_00842_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[118][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12342_ (.D(_00843_),
    .CLK(net346),
    .Q(\u_cpu.rf_ram.memory[118][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12343_ (.D(_00844_),
    .CLK(net346),
    .Q(\u_cpu.rf_ram.memory[118][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12344_ (.D(_00845_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[118][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12345_ (.D(_00846_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[118][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12346_ (.D(_00847_),
    .CLK(net455),
    .Q(\u_cpu.rf_ram.memory[118][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12347_ (.D(_00848_),
    .CLK(net452),
    .Q(\u_cpu.rf_ram.memory[118][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12348_ (.D(_00849_),
    .CLK(net452),
    .Q(\u_cpu.rf_ram.memory[118][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12349_ (.D(_00850_),
    .CLK(net472),
    .Q(\u_cpu.rf_ram.memory[121][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12350_ (.D(_00851_),
    .CLK(net361),
    .Q(\u_cpu.rf_ram.memory[121][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12351_ (.D(_00852_),
    .CLK(net364),
    .Q(\u_cpu.rf_ram.memory[121][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12352_ (.D(_00853_),
    .CLK(net364),
    .Q(\u_cpu.rf_ram.memory[121][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12353_ (.D(_00854_),
    .CLK(net364),
    .Q(\u_cpu.rf_ram.memory[121][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12354_ (.D(_00855_),
    .CLK(net362),
    .Q(\u_cpu.rf_ram.memory[121][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12355_ (.D(_00856_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[121][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12356_ (.D(_00857_),
    .CLK(net472),
    .Q(\u_cpu.rf_ram.memory[121][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12357_ (.D(_00858_),
    .CLK(net423),
    .Q(\u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12358_ (.D(_00859_),
    .CLK(net423),
    .Q(\u_cpu.rf_ram.memory[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12359_ (.D(_00860_),
    .CLK(net441),
    .Q(\u_cpu.rf_ram.memory[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12360_ (.D(_00861_),
    .CLK(net441),
    .Q(\u_cpu.rf_ram.memory[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12361_ (.D(_00862_),
    .CLK(net423),
    .Q(\u_cpu.rf_ram.memory[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12362_ (.D(_00863_),
    .CLK(net423),
    .Q(\u_cpu.rf_ram.memory[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12363_ (.D(_00864_),
    .CLK(net414),
    .Q(\u_cpu.rf_ram.memory[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12364_ (.D(_00865_),
    .CLK(net414),
    .Q(\u_cpu.rf_ram.memory[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12365_ (.D(_00866_),
    .CLK(net422),
    .Q(\u_cpu.rf_ram.memory[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12366_ (.D(_00867_),
    .CLK(net422),
    .Q(\u_cpu.rf_ram.memory[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12367_ (.D(_00868_),
    .CLK(net422),
    .Q(\u_cpu.rf_ram.memory[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12368_ (.D(_00869_),
    .CLK(net422),
    .Q(\u_cpu.rf_ram.memory[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12369_ (.D(_00870_),
    .CLK(net422),
    .Q(\u_cpu.rf_ram.memory[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12370_ (.D(_00871_),
    .CLK(net423),
    .Q(\u_cpu.rf_ram.memory[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12371_ (.D(_00872_),
    .CLK(net414),
    .Q(\u_cpu.rf_ram.memory[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12372_ (.D(_00873_),
    .CLK(net417),
    .Q(\u_cpu.rf_ram.memory[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12373_ (.D(_00874_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[112][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12374_ (.D(_00875_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[112][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12375_ (.D(_00876_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[112][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12376_ (.D(_00877_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[112][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12377_ (.D(_00878_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[112][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12378_ (.D(_00879_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[112][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12379_ (.D(_00880_),
    .CLK(net478),
    .Q(\u_cpu.rf_ram.memory[112][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12380_ (.D(_00881_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[112][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12381_ (.D(_00882_),
    .CLK(net472),
    .Q(\u_cpu.rf_ram.memory[122][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12382_ (.D(_00883_),
    .CLK(net472),
    .Q(\u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12383_ (.D(_00884_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[122][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12384_ (.D(_00885_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[122][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12385_ (.D(_00886_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[122][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12386_ (.D(_00887_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[122][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12387_ (.D(_00888_),
    .CLK(net473),
    .Q(\u_cpu.rf_ram.memory[122][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12388_ (.D(_00889_),
    .CLK(net472),
    .Q(\u_cpu.rf_ram.memory[122][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12389_ (.D(_00890_),
    .CLK(net474),
    .Q(\u_cpu.rf_ram.memory[115][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12390_ (.D(_00891_),
    .CLK(net475),
    .Q(\u_cpu.rf_ram.memory[115][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12391_ (.D(_00892_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[115][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12392_ (.D(_00893_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[115][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12393_ (.D(_00894_),
    .CLK(net482),
    .Q(\u_cpu.rf_ram.memory[115][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12394_ (.D(_00895_),
    .CLK(net491),
    .Q(\u_cpu.rf_ram.memory[115][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12395_ (.D(_00896_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[115][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12396_ (.D(_00897_),
    .CLK(net474),
    .Q(\u_cpu.rf_ram.memory[115][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12397_ (.D(_00898_),
    .CLK(net458),
    .Q(\u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12398_ (.D(_00899_),
    .CLK(net458),
    .Q(\u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12399_ (.D(_00900_),
    .CLK(net454),
    .Q(\u_cpu.rf_ram.memory[116][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12400_ (.D(_00901_),
    .CLK(net459),
    .Q(\u_cpu.rf_ram.memory[116][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12401_ (.D(_00902_),
    .CLK(net455),
    .Q(\u_cpu.rf_ram.memory[116][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12402_ (.D(_00903_),
    .CLK(net455),
    .Q(\u_cpu.rf_ram.memory[116][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12403_ (.D(_00904_),
    .CLK(net455),
    .Q(\u_cpu.rf_ram.memory[116][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12404_ (.D(_00905_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[116][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12405_ (.D(_00906_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[33][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12406_ (.D(_00907_),
    .CLK(net465),
    .Q(\u_cpu.rf_ram.memory[33][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12407_ (.D(_00908_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[33][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12408_ (.D(_00909_),
    .CLK(net486),
    .Q(\u_cpu.rf_ram.memory[33][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12409_ (.D(_00910_),
    .CLK(net486),
    .Q(\u_cpu.rf_ram.memory[33][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12410_ (.D(_00911_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[33][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12411_ (.D(_00912_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12412_ (.D(_00913_),
    .CLK(net465),
    .Q(\u_cpu.rf_ram.memory[33][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12413_ (.D(_00914_),
    .CLK(net247),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12414_ (.D(_00915_),
    .CLK(net249),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12415_ (.D(_00916_),
    .CLK(net249),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12416_ (.D(_00917_),
    .CLK(net247),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12417_ (.D(_00918_),
    .CLK(net247),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12418_ (.D(_00919_),
    .CLK(net248),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12419_ (.D(_00920_),
    .CLK(net248),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12420_ (.D(_00921_),
    .CLK(net235),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12421_ (.D(_00922_),
    .CLK(net235),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12422_ (.D(_00923_),
    .CLK(net234),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12423_ (.D(_00924_),
    .CLK(net234),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12424_ (.D(_00925_),
    .CLK(net233),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12425_ (.D(_00926_),
    .CLK(net233),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12426_ (.D(_00927_),
    .CLK(net49),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12427_ (.D(_00928_),
    .CLK(net47),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12428_ (.D(_00929_),
    .CLK(net47),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12429_ (.D(_00930_),
    .CLK(net49),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12430_ (.D(_00931_),
    .CLK(net49),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12431_ (.D(_00932_),
    .CLK(net233),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12432_ (.D(_00933_),
    .CLK(net233),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12433_ (.D(_00934_),
    .CLK(net233),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12434_ (.D(_00935_),
    .CLK(net235),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12435_ (.D(_00936_),
    .CLK(net236),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12436_ (.D(_00937_),
    .CLK(net246),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12437_ (.D(_00938_),
    .CLK(net246),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12438_ (.D(_00939_),
    .CLK(net246),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12439_ (.D(_00940_),
    .CLK(net246),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12440_ (.D(_00941_),
    .CLK(net246),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12441_ (.D(_00942_),
    .CLK(net247),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12442_ (.D(_00943_),
    .CLK(net249),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12443_ (.D(_00944_),
    .CLK(net249),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12444_ (.D(_00945_),
    .CLK(net249),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12445_ (.D(_00946_),
    .CLK(net474),
    .Q(\u_cpu.rf_ram.memory[113][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12446_ (.D(_00947_),
    .CLK(net475),
    .Q(\u_cpu.rf_ram.memory[113][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12447_ (.D(_00948_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[113][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12448_ (.D(_00949_),
    .CLK(net478),
    .Q(\u_cpu.rf_ram.memory[113][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12449_ (.D(_00950_),
    .CLK(net482),
    .Q(\u_cpu.rf_ram.memory[113][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12450_ (.D(_00951_),
    .CLK(net482),
    .Q(\u_cpu.rf_ram.memory[113][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12451_ (.D(_00952_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[113][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12452_ (.D(_00953_),
    .CLK(net474),
    .Q(\u_cpu.rf_ram.memory[113][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12453_ (.D(_00954_),
    .CLK(net252),
    .Q(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12454_ (.D(_00955_),
    .CLK(net252),
    .Q(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12455_ (.D(_00956_),
    .CLK(net252),
    .Q(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12456_ (.D(_00957_),
    .CLK(net253),
    .Q(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12457_ (.D(_00958_),
    .CLK(net252),
    .Q(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12458_ (.D(_00959_),
    .CLK(net253),
    .Q(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12459_ (.D(_00960_),
    .CLK(net254),
    .Q(\u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12460_ (.D(_00961_),
    .CLK(net253),
    .Q(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12461_ (.D(_00962_),
    .CLK(net253),
    .Q(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12462_ (.D(_00963_),
    .CLK(net253),
    .Q(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12463_ (.D(_00964_),
    .CLK(net263),
    .Q(\u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12464_ (.D(_00965_),
    .CLK(net474),
    .Q(\u_cpu.rf_ram.memory[114][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12465_ (.D(_00966_),
    .CLK(net486),
    .Q(\u_cpu.rf_ram.memory[114][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12466_ (.D(_00967_),
    .CLK(net490),
    .Q(\u_cpu.rf_ram.memory[114][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12467_ (.D(_00968_),
    .CLK(net491),
    .Q(\u_cpu.rf_ram.memory[114][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12468_ (.D(_00969_),
    .CLK(net491),
    .Q(\u_cpu.rf_ram.memory[114][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12469_ (.D(_00970_),
    .CLK(net491),
    .Q(\u_cpu.rf_ram.memory[114][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12470_ (.D(_00971_),
    .CLK(net490),
    .Q(\u_cpu.rf_ram.memory[114][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12471_ (.D(_00972_),
    .CLK(net475),
    .Q(\u_cpu.rf_ram.memory[114][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12472_ (.D(_00973_),
    .CLK(net279),
    .Q(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12473_ (.D(_00974_),
    .CLK(net237),
    .Q(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12474_ (.D(_00975_),
    .CLK(net259),
    .Q(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12475_ (.D(_00976_),
    .CLK(net237),
    .Q(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12476_ (.D(_00977_),
    .CLK(net238),
    .Q(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12477_ (.D(_00978_),
    .CLK(net238),
    .Q(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12478_ (.D(_00979_),
    .CLK(net240),
    .Q(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12479_ (.D(_00980_),
    .CLK(net240),
    .Q(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12480_ (.D(_00981_),
    .CLK(net240),
    .Q(\u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12481_ (.D(_00982_),
    .CLK(net240),
    .Q(\u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12482_ (.D(_00983_),
    .CLK(net239),
    .Q(\u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12483_ (.D(_00984_),
    .CLK(net241),
    .Q(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12484_ (.D(_00985_),
    .CLK(net242),
    .Q(\u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12485_ (.D(_00986_),
    .CLK(net243),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12486_ (.D(_00987_),
    .CLK(net242),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12487_ (.D(_00988_),
    .CLK(net242),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12488_ (.D(_00989_),
    .CLK(net242),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12489_ (.D(_00990_),
    .CLK(net242),
    .Q(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12490_ (.D(_00991_),
    .CLK(net237),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12491_ (.D(_00992_),
    .CLK(net237),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12492_ (.D(_00993_),
    .CLK(net237),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12493_ (.D(_00994_),
    .CLK(net53),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12494_ (.D(_00995_),
    .CLK(net240),
    .Q(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12495_ (.D(_00996_),
    .CLK(net316),
    .Q(\u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12496_ (.D(_00997_),
    .CLK(net492),
    .Q(\u_cpu.rf_ram.memory[32][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12497_ (.D(_00998_),
    .CLK(net492),
    .Q(\u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12498_ (.D(_00999_),
    .CLK(net492),
    .Q(\u_cpu.rf_ram.memory[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12499_ (.D(_01000_),
    .CLK(net493),
    .Q(\u_cpu.rf_ram.memory[32][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12500_ (.D(_01001_),
    .CLK(net491),
    .Q(\u_cpu.rf_ram.memory[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12501_ (.D(_01002_),
    .CLK(net490),
    .Q(\u_cpu.rf_ram.memory[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12502_ (.D(_01003_),
    .CLK(net490),
    .Q(\u_cpu.rf_ram.memory[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12503_ (.D(_01004_),
    .CLK(net490),
    .Q(\u_cpu.rf_ram.memory[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12504_ (.D(_01005_),
    .CLK(net186),
    .Q(\u_cpu.rf_ram.memory[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12505_ (.D(_01006_),
    .CLK(net186),
    .Q(\u_cpu.rf_ram.memory[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12506_ (.D(_01007_),
    .CLK(net172),
    .Q(\u_cpu.rf_ram.memory[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12507_ (.D(_01008_),
    .CLK(net176),
    .Q(\u_cpu.rf_ram.memory[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12508_ (.D(_01009_),
    .CLK(net172),
    .Q(\u_cpu.rf_ram.memory[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12509_ (.D(_01010_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12510_ (.D(_01011_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12511_ (.D(_01012_),
    .CLK(net183),
    .Q(\u_cpu.rf_ram.memory[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12512_ (.D(_01013_),
    .CLK(net255),
    .Q(\u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12513_ (.D(_01014_),
    .CLK(net307),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12514_ (.D(_01015_),
    .CLK(net307),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12515_ (.D(_01016_),
    .CLK(net307),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12516_ (.D(_01017_),
    .CLK(net307),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12517_ (.D(_01018_),
    .CLK(net307),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12518_ (.D(_01019_),
    .CLK(net311),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12519_ (.D(_01020_),
    .CLK(net311),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12520_ (.D(_01021_),
    .CLK(net311),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12521_ (.D(_01022_),
    .CLK(net322),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12522_ (.D(_01023_),
    .CLK(net311),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12523_ (.D(_01024_),
    .CLK(net322),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12524_ (.D(_01025_),
    .CLK(net322),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12525_ (.D(_01026_),
    .CLK(net322),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12526_ (.D(_01027_),
    .CLK(net322),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12527_ (.D(_01028_),
    .CLK(net324),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12528_ (.D(_01029_),
    .CLK(net324),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12529_ (.D(_01030_),
    .CLK(net324),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12530_ (.D(_01031_),
    .CLK(net324),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12531_ (.D(_01032_),
    .CLK(net324),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12532_ (.D(_01033_),
    .CLK(net325),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12533_ (.D(_01034_),
    .CLK(net329),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12534_ (.D(_01035_),
    .CLK(net330),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12535_ (.D(_01036_),
    .CLK(net330),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12536_ (.D(_01037_),
    .CLK(net330),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12537_ (.D(_01038_),
    .CLK(net328),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12538_ (.D(_01039_),
    .CLK(net328),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12539_ (.D(_01040_),
    .CLK(net328),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12540_ (.D(_01041_),
    .CLK(net318),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12541_ (.D(_01042_),
    .CLK(net318),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12542_ (.D(_01043_),
    .CLK(net318),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12543_ (.D(_00022_),
    .CLK(net252),
    .Q(\u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12544_ (.D(_01044_),
    .CLK(net255),
    .Q(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12545_ (.D(_01045_),
    .CLK(net254),
    .Q(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12546_ (.D(_01046_),
    .CLK(net187),
    .Q(\u_cpu.rf_ram.memory[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12547_ (.D(_01047_),
    .CLK(net187),
    .Q(\u_cpu.rf_ram.memory[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12548_ (.D(_01048_),
    .CLK(net172),
    .Q(\u_cpu.rf_ram.memory[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12549_ (.D(_01049_),
    .CLK(net173),
    .Q(\u_cpu.rf_ram.memory[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12550_ (.D(_01050_),
    .CLK(net173),
    .Q(\u_cpu.rf_ram.memory[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12551_ (.D(_01051_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12552_ (.D(_01052_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12553_ (.D(_01053_),
    .CLK(net184),
    .Q(\u_cpu.rf_ram.memory[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12554_ (.D(_00024_),
    .CLK(net313),
    .Q(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12555_ (.D(_00023_),
    .CLK(net313),
    .Q(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12556_ (.D(_01054_),
    .CLK(net313),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12557_ (.D(_01055_),
    .CLK(net250),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12558_ (.D(_01056_),
    .CLK(net250),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12559_ (.D(_01057_),
    .CLK(net308),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12560_ (.D(_01058_),
    .CLK(net308),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12561_ (.D(_01059_),
    .CLK(net309),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12562_ (.D(_01060_),
    .CLK(net309),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12563_ (.D(_01061_),
    .CLK(net309),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12564_ (.D(_01062_),
    .CLK(net309),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12565_ (.D(_01063_),
    .CLK(net309),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12566_ (.D(_01064_),
    .CLK(net310),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12567_ (.D(_01065_),
    .CLK(net310),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12568_ (.D(_01066_),
    .CLK(net323),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12569_ (.D(_01067_),
    .CLK(net323),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12570_ (.D(_01068_),
    .CLK(net323),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12571_ (.D(_01069_),
    .CLK(net327),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12572_ (.D(_01070_),
    .CLK(net323),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12573_ (.D(_01071_),
    .CLK(net325),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12574_ (.D(_01072_),
    .CLK(net325),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12575_ (.D(_01073_),
    .CLK(net325),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12576_ (.D(_01074_),
    .CLK(net329),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12577_ (.D(_01075_),
    .CLK(net329),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12578_ (.D(_01076_),
    .CLK(net329),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12579_ (.D(_01077_),
    .CLK(net330),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12580_ (.D(_01078_),
    .CLK(net329),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12581_ (.D(_01079_),
    .CLK(net327),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12582_ (.D(_01080_),
    .CLK(net327),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12583_ (.D(_01081_),
    .CLK(net327),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12584_ (.D(_01082_),
    .CLK(net327),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12585_ (.D(_01083_),
    .CLK(net319),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12586_ (.D(_01084_),
    .CLK(net319),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12587_ (.D(_01085_),
    .CLK(net319),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12588_ (.D(_01086_),
    .CLK(net172),
    .Q(\u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12589_ (.D(_01087_),
    .CLK(net172),
    .Q(\u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12590_ (.D(_01088_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[109][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12591_ (.D(_01089_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[109][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12592_ (.D(_01090_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[109][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12593_ (.D(_01091_),
    .CLK(net171),
    .Q(\u_cpu.rf_ram.memory[109][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12594_ (.D(_01092_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[109][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12595_ (.D(_01093_),
    .CLK(net166),
    .Q(\u_cpu.rf_ram.memory[109][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12596_ (.D(_00021_),
    .CLK(net280),
    .Q(\u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12597_ (.D(_01094_),
    .CLK(net441),
    .Q(\u_cpu.rf_ram.memory[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12598_ (.D(_01095_),
    .CLK(net441),
    .Q(\u_cpu.rf_ram.memory[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12599_ (.D(_01096_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12600_ (.D(_01097_),
    .CLK(net446),
    .Q(\u_cpu.rf_ram.memory[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12601_ (.D(_01098_),
    .CLK(net446),
    .Q(\u_cpu.rf_ram.memory[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12602_ (.D(_01099_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12603_ (.D(_01100_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12604_ (.D(_01101_),
    .CLK(net442),
    .Q(\u_cpu.rf_ram.memory[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12605_ (.D(_01102_),
    .CLK(net443),
    .Q(\u_cpu.rf_ram.memory[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12606_ (.D(_01103_),
    .CLK(net443),
    .Q(\u_cpu.rf_ram.memory[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12607_ (.D(_01104_),
    .CLK(net447),
    .Q(\u_cpu.rf_ram.memory[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12608_ (.D(_01105_),
    .CLK(net447),
    .Q(\u_cpu.rf_ram.memory[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12609_ (.D(_01106_),
    .CLK(net447),
    .Q(\u_cpu.rf_ram.memory[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12610_ (.D(_01107_),
    .CLK(net443),
    .Q(\u_cpu.rf_ram.memory[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12611_ (.D(_01108_),
    .CLK(net444),
    .Q(\u_cpu.rf_ram.memory[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12612_ (.D(_01109_),
    .CLK(net444),
    .Q(\u_cpu.rf_ram.memory[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12613_ (.D(_01110_),
    .CLK(net151),
    .Q(\u_cpu.rf_ram.memory[93][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12614_ (.D(_01111_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[93][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12615_ (.D(_01112_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[93][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12616_ (.D(_01113_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[93][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12617_ (.D(_01114_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[93][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12618_ (.D(_01115_),
    .CLK(net146),
    .Q(\u_cpu.rf_ram.memory[93][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12619_ (.D(_01116_),
    .CLK(net146),
    .Q(\u_cpu.rf_ram.memory[93][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12620_ (.D(_01117_),
    .CLK(net148),
    .Q(\u_cpu.rf_ram.memory[93][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12621_ (.D(_01118_),
    .CLK(net263),
    .Q(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12622_ (.D(_01119_),
    .CLK(net263),
    .Q(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12623_ (.D(_01120_),
    .CLK(net263),
    .Q(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12624_ (.D(_01121_),
    .CLK(net263),
    .Q(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12625_ (.D(_01122_),
    .CLK(net266),
    .Q(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12626_ (.D(_01123_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[97][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12627_ (.D(_01124_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[97][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12628_ (.D(_01125_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[97][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12629_ (.D(_01126_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[97][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12630_ (.D(_01127_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[97][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12631_ (.D(_01128_),
    .CLK(net156),
    .Q(\u_cpu.rf_ram.memory[97][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12632_ (.D(_01129_),
    .CLK(net154),
    .Q(\u_cpu.rf_ram.memory[97][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12633_ (.D(_01130_),
    .CLK(net194),
    .Q(\u_cpu.rf_ram.memory[97][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12634_ (.D(_01131_),
    .CLK(net151),
    .Q(\u_cpu.rf_ram.memory[94][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12635_ (.D(_01132_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[94][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12636_ (.D(_01133_),
    .CLK(net146),
    .Q(\u_cpu.rf_ram.memory[94][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12637_ (.D(_01134_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[94][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12638_ (.D(_01135_),
    .CLK(net146),
    .Q(\u_cpu.rf_ram.memory[94][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12639_ (.D(_01136_),
    .CLK(net145),
    .Q(\u_cpu.rf_ram.memory[94][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12640_ (.D(_01137_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[94][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12641_ (.D(_01138_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[94][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12642_ (.D(_01139_),
    .CLK(net148),
    .Q(\u_cpu.rf_ram.memory[95][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12643_ (.D(_01140_),
    .CLK(net147),
    .Q(\u_cpu.rf_ram.memory[95][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12644_ (.D(_01141_),
    .CLK(net147),
    .Q(\u_cpu.rf_ram.memory[95][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12645_ (.D(_01142_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[95][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12646_ (.D(_01143_),
    .CLK(net146),
    .Q(\u_cpu.rf_ram.memory[95][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12647_ (.D(_01144_),
    .CLK(net145),
    .Q(\u_cpu.rf_ram.memory[95][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12648_ (.D(_01145_),
    .CLK(net144),
    .Q(\u_cpu.rf_ram.memory[95][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12649_ (.D(_01146_),
    .CLK(net144),
    .Q(\u_cpu.rf_ram.memory[95][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12650_ (.D(_01147_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[96][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12651_ (.D(_01148_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[96][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12652_ (.D(_01149_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[96][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12653_ (.D(_01150_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[96][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12654_ (.D(_01151_),
    .CLK(net160),
    .Q(\u_cpu.rf_ram.memory[96][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12655_ (.D(_01152_),
    .CLK(net156),
    .Q(\u_cpu.rf_ram.memory[96][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12656_ (.D(_01153_),
    .CLK(net154),
    .Q(\u_cpu.rf_ram.memory[96][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12657_ (.D(_01154_),
    .CLK(net194),
    .Q(\u_cpu.rf_ram.memory[96][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12658_ (.D(_01155_),
    .CLK(net241),
    .Q(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12659_ (.D(_01156_),
    .CLK(net236),
    .Q(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12660_ (.D(_01157_),
    .CLK(net176),
    .Q(\u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12661_ (.D(_01158_),
    .CLK(net176),
    .Q(\u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12662_ (.D(_01159_),
    .CLK(net197),
    .Q(\u_cpu.rf_ram.memory[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12663_ (.D(_01160_),
    .CLK(net197),
    .Q(\u_cpu.rf_ram.memory[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12664_ (.D(_01161_),
    .CLK(net197),
    .Q(\u_cpu.rf_ram.memory[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12665_ (.D(_01162_),
    .CLK(net177),
    .Q(\u_cpu.rf_ram.memory[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12666_ (.D(_01163_),
    .CLK(net177),
    .Q(\u_cpu.rf_ram.memory[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12667_ (.D(_01164_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12668_ (.D(_01165_),
    .CLK(net47),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12669_ (.D(_01166_),
    .CLK(net47),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12670_ (.D(_01167_),
    .CLK(net48),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12671_ (.D(_01168_),
    .CLK(net49),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12672_ (.D(_01169_),
    .CLK(net49),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12673_ (.D(_01170_),
    .CLK(net50),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12674_ (.D(_01171_),
    .CLK(net50),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12675_ (.D(_01172_),
    .CLK(net48),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12676_ (.D(_01173_),
    .CLK(net48),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12677_ (.D(_01174_),
    .CLK(net234),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12678_ (.D(_01175_),
    .CLK(net50),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12679_ (.D(_01176_),
    .CLK(net47),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12680_ (.D(_01177_),
    .CLK(net46),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12681_ (.D(_01178_),
    .CLK(net46),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12682_ (.D(_01179_),
    .CLK(net46),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12683_ (.D(_01180_),
    .CLK(net46),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12684_ (.D(_01181_),
    .CLK(net170),
    .Q(\u_cpu.rf_ram.memory[101][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12685_ (.D(_01182_),
    .CLK(net170),
    .Q(\u_cpu.rf_ram.memory[101][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12686_ (.D(_01183_),
    .CLK(net194),
    .Q(\u_cpu.rf_ram.memory[101][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12687_ (.D(_01184_),
    .CLK(net194),
    .Q(\u_cpu.rf_ram.memory[101][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12688_ (.D(_01185_),
    .CLK(net194),
    .Q(\u_cpu.rf_ram.memory[101][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12689_ (.D(_01186_),
    .CLK(net170),
    .Q(\u_cpu.rf_ram.memory[101][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12690_ (.D(_01187_),
    .CLK(net170),
    .Q(\u_cpu.rf_ram.memory[101][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12691_ (.D(_01188_),
    .CLK(net170),
    .Q(\u_cpu.rf_ram.memory[101][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12692_ (.D(_01189_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12693_ (.D(_01190_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12694_ (.D(_01191_),
    .CLK(net153),
    .Q(\u_cpu.rf_ram.memory[102][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12695_ (.D(_01192_),
    .CLK(net153),
    .Q(\u_cpu.rf_ram.memory[102][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12696_ (.D(_01193_),
    .CLK(net153),
    .Q(\u_cpu.rf_ram.memory[102][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12697_ (.D(_01194_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[102][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12698_ (.D(_01195_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[102][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12699_ (.D(_01196_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[102][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12700_ (.D(_01197_),
    .CLK(net137),
    .Q(\u_cpu.rf_ram.memory[103][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12701_ (.D(_01198_),
    .CLK(net137),
    .Q(\u_cpu.rf_ram.memory[103][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12702_ (.D(_01199_),
    .CLK(net154),
    .Q(\u_cpu.rf_ram.memory[103][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12703_ (.D(_01200_),
    .CLK(net154),
    .Q(\u_cpu.rf_ram.memory[103][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12704_ (.D(_01201_),
    .CLK(net154),
    .Q(\u_cpu.rf_ram.memory[103][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12705_ (.D(_01202_),
    .CLK(net137),
    .Q(\u_cpu.rf_ram.memory[103][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12706_ (.D(_01203_),
    .CLK(net137),
    .Q(\u_cpu.rf_ram.memory[103][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12707_ (.D(_01204_),
    .CLK(net171),
    .Q(\u_cpu.rf_ram.memory[103][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12708_ (.D(_01205_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12709_ (.D(_01206_),
    .CLK(net135),
    .Q(\u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12710_ (.D(_01207_),
    .CLK(net151),
    .Q(\u_cpu.rf_ram.memory[104][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12711_ (.D(_01208_),
    .CLK(net151),
    .Q(\u_cpu.rf_ram.memory[104][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12712_ (.D(_01209_),
    .CLK(net151),
    .Q(\u_cpu.rf_ram.memory[104][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12713_ (.D(_01210_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[104][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12714_ (.D(_01211_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[104][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12715_ (.D(_01212_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[104][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12716_ (.D(_01213_),
    .CLK(net155),
    .Q(\u_cpu.rf_ram.memory[99][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12717_ (.D(_01214_),
    .CLK(net155),
    .Q(\u_cpu.rf_ram.memory[99][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12718_ (.D(_01215_),
    .CLK(net155),
    .Q(\u_cpu.rf_ram.memory[99][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12719_ (.D(_01216_),
    .CLK(net155),
    .Q(\u_cpu.rf_ram.memory[99][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12720_ (.D(_01217_),
    .CLK(net156),
    .Q(\u_cpu.rf_ram.memory[99][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12721_ (.D(_01218_),
    .CLK(net155),
    .Q(\u_cpu.rf_ram.memory[99][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12722_ (.D(_01219_),
    .CLK(net153),
    .Q(\u_cpu.rf_ram.memory[99][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12723_ (.D(_01220_),
    .CLK(net153),
    .Q(\u_cpu.rf_ram.memory[99][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12724_ (.D(_01221_),
    .CLK(net124),
    .Q(\u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12725_ (.D(_01222_),
    .CLK(net124),
    .Q(\u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12726_ (.D(_01223_),
    .CLK(net128),
    .Q(\u_cpu.rf_ram.memory[79][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12727_ (.D(_01224_),
    .CLK(net128),
    .Q(\u_cpu.rf_ram.memory[79][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12728_ (.D(_01225_),
    .CLK(net128),
    .Q(\u_cpu.rf_ram.memory[79][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12729_ (.D(_01226_),
    .CLK(net124),
    .Q(\u_cpu.rf_ram.memory[79][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12730_ (.D(_01227_),
    .CLK(net124),
    .Q(\u_cpu.rf_ram.memory[79][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12731_ (.D(_01228_),
    .CLK(net124),
    .Q(\u_cpu.rf_ram.memory[79][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12732_ (.D(_01229_),
    .CLK(net120),
    .Q(\u_cpu.rf_ram.memory[105][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12733_ (.D(_01230_),
    .CLK(net120),
    .Q(\u_cpu.rf_ram.memory[105][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12734_ (.D(_01231_),
    .CLK(net148),
    .Q(\u_cpu.rf_ram.memory[105][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12735_ (.D(_01232_),
    .CLK(net148),
    .Q(\u_cpu.rf_ram.memory[105][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12736_ (.D(_01233_),
    .CLK(net148),
    .Q(\u_cpu.rf_ram.memory[105][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12737_ (.D(_01234_),
    .CLK(net120),
    .Q(\u_cpu.rf_ram.memory[105][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12738_ (.D(_01235_),
    .CLK(net121),
    .Q(\u_cpu.rf_ram.memory[105][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12739_ (.D(_01236_),
    .CLK(net121),
    .Q(\u_cpu.rf_ram.memory[105][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12740_ (.D(_01237_),
    .CLK(net115),
    .Q(\u_cpu.rf_ram.memory[106][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12741_ (.D(_01238_),
    .CLK(net115),
    .Q(\u_cpu.rf_ram.memory[106][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12742_ (.D(_01239_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[106][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12743_ (.D(_01240_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[106][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12744_ (.D(_01241_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[106][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12745_ (.D(_01242_),
    .CLK(net115),
    .Q(\u_cpu.rf_ram.memory[106][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12746_ (.D(_01243_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[106][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12747_ (.D(_01244_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[106][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12748_ (.D(_01245_),
    .CLK(net115),
    .Q(\u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12749_ (.D(_01246_),
    .CLK(net115),
    .Q(\u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12750_ (.D(_01247_),
    .CLK(net144),
    .Q(\u_cpu.rf_ram.memory[107][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12751_ (.D(_01248_),
    .CLK(net144),
    .Q(\u_cpu.rf_ram.memory[107][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12752_ (.D(_01249_),
    .CLK(net145),
    .Q(\u_cpu.rf_ram.memory[107][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12753_ (.D(_01250_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[107][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12754_ (.D(_01251_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[107][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12755_ (.D(_01252_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[107][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12756_ (.D(_01253_),
    .CLK(net186),
    .Q(\u_cpu.rf_ram.memory[83][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12757_ (.D(_01254_),
    .CLK(net186),
    .Q(\u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12758_ (.D(_01255_),
    .CLK(net207),
    .Q(\u_cpu.rf_ram.memory[83][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12759_ (.D(_01256_),
    .CLK(net207),
    .Q(\u_cpu.rf_ram.memory[83][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12760_ (.D(_01257_),
    .CLK(net208),
    .Q(\u_cpu.rf_ram.memory[83][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12761_ (.D(_01258_),
    .CLK(net207),
    .Q(\u_cpu.rf_ram.memory[83][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12762_ (.D(_01259_),
    .CLK(net207),
    .Q(\u_cpu.rf_ram.memory[83][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12763_ (.D(_01260_),
    .CLK(net186),
    .Q(\u_cpu.rf_ram.memory[83][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12764_ (.D(_01261_),
    .CLK(net171),
    .Q(\u_cpu.rf_ram.memory[108][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12765_ (.D(_01262_),
    .CLK(net171),
    .Q(\u_cpu.rf_ram.memory[108][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12766_ (.D(_01263_),
    .CLK(net138),
    .Q(\u_cpu.rf_ram.memory[108][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12767_ (.D(_01264_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[108][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12768_ (.D(_01265_),
    .CLK(net138),
    .Q(\u_cpu.rf_ram.memory[108][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12769_ (.D(_01266_),
    .CLK(net138),
    .Q(\u_cpu.rf_ram.memory[108][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12770_ (.D(_01267_),
    .CLK(net138),
    .Q(\u_cpu.rf_ram.memory[108][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12771_ (.D(_01268_),
    .CLK(net129),
    .Q(\u_cpu.rf_ram.memory[108][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12772_ (.D(_01269_),
    .CLK(net12),
    .Q(\u_cpu.rf_ram.memory[69][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12773_ (.D(_01270_),
    .CLK(net12),
    .Q(\u_cpu.rf_ram.memory[69][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12774_ (.D(_01271_),
    .CLK(net11),
    .Q(\u_cpu.rf_ram.memory[69][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12775_ (.D(_01272_),
    .CLK(net11),
    .Q(\u_cpu.rf_ram.memory[69][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12776_ (.D(_01273_),
    .CLK(net13),
    .Q(\u_cpu.rf_ram.memory[69][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12777_ (.D(_01274_),
    .CLK(net12),
    .Q(\u_cpu.rf_ram.memory[69][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12778_ (.D(_01275_),
    .CLK(net13),
    .Q(\u_cpu.rf_ram.memory[69][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12779_ (.D(_01276_),
    .CLK(net18),
    .Q(\u_cpu.rf_ram.memory[69][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12780_ (.D(_01277_),
    .CLK(net102),
    .Q(\u_cpu.rf_ram.memory[84][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12781_ (.D(_01278_),
    .CLK(net102),
    .Q(\u_cpu.rf_ram.memory[84][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12782_ (.D(_01279_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[84][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12783_ (.D(_01280_),
    .CLK(net118),
    .Q(\u_cpu.rf_ram.memory[84][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12784_ (.D(_01281_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[84][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12785_ (.D(_01282_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[84][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12786_ (.D(_01283_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[84][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12787_ (.D(_01284_),
    .CLK(net108),
    .Q(\u_cpu.rf_ram.memory[84][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12788_ (.D(_01285_),
    .CLK(net70),
    .Q(\u_cpu.rf_ram.memory[59][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12789_ (.D(_01286_),
    .CLK(net70),
    .Q(\u_cpu.rf_ram.memory[59][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12790_ (.D(_01287_),
    .CLK(net73),
    .Q(\u_cpu.rf_ram.memory[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12791_ (.D(_01288_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[59][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12792_ (.D(_01289_),
    .CLK(net70),
    .Q(\u_cpu.rf_ram.memory[59][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12793_ (.D(_01290_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12794_ (.D(_01291_),
    .CLK(net39),
    .Q(\u_cpu.rf_ram.memory[59][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12795_ (.D(_01292_),
    .CLK(net39),
    .Q(\u_cpu.rf_ram.memory[59][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12796_ (.D(_01293_),
    .CLK(net412),
    .Q(\u_cpu.rf_ram.memory[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12797_ (.D(_01294_),
    .CLK(net412),
    .Q(\u_cpu.rf_ram.memory[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12798_ (.D(_01295_),
    .CLK(net412),
    .Q(\u_cpu.rf_ram.memory[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12799_ (.D(_01296_),
    .CLK(net413),
    .Q(\u_cpu.rf_ram.memory[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12800_ (.D(_01297_),
    .CLK(net413),
    .Q(\u_cpu.rf_ram.memory[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12801_ (.D(_01298_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12802_ (.D(_01299_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12803_ (.D(_01300_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12804_ (.D(_01301_),
    .CLK(net100),
    .Q(\u_cpu.rf_ram.memory[85][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12805_ (.D(_01302_),
    .CLK(net103),
    .Q(\u_cpu.rf_ram.memory[85][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12806_ (.D(_01303_),
    .CLK(net111),
    .Q(\u_cpu.rf_ram.memory[85][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12807_ (.D(_01304_),
    .CLK(net119),
    .Q(\u_cpu.rf_ram.memory[85][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12808_ (.D(_01305_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[85][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12809_ (.D(_01306_),
    .CLK(net111),
    .Q(\u_cpu.rf_ram.memory[85][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12810_ (.D(_01307_),
    .CLK(net119),
    .Q(\u_cpu.rf_ram.memory[85][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12811_ (.D(_01308_),
    .CLK(net108),
    .Q(\u_cpu.rf_ram.memory[85][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12812_ (.D(_01309_),
    .CLK(net125),
    .Q(\u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12813_ (.D(_01310_),
    .CLK(net131),
    .Q(\u_cpu.rf_ram.memory[110][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12814_ (.D(_01311_),
    .CLK(net131),
    .Q(\u_cpu.rf_ram.memory[110][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12815_ (.D(_01312_),
    .CLK(net131),
    .Q(\u_cpu.rf_ram.memory[110][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12816_ (.D(_01313_),
    .CLK(net132),
    .Q(\u_cpu.rf_ram.memory[110][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12817_ (.D(_01314_),
    .CLK(net131),
    .Q(\u_cpu.rf_ram.memory[110][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12818_ (.D(_01315_),
    .CLK(net131),
    .Q(\u_cpu.rf_ram.memory[110][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12819_ (.D(_01316_),
    .CLK(net125),
    .Q(\u_cpu.rf_ram.memory[110][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12820_ (.D(_01317_),
    .CLK(net100),
    .Q(\u_cpu.rf_ram.memory[86][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12821_ (.D(_01318_),
    .CLK(net101),
    .Q(\u_cpu.rf_ram.memory[86][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12822_ (.D(_01319_),
    .CLK(net111),
    .Q(\u_cpu.rf_ram.memory[86][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12823_ (.D(_01320_),
    .CLK(net118),
    .Q(\u_cpu.rf_ram.memory[86][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12824_ (.D(_01321_),
    .CLK(net113),
    .Q(\u_cpu.rf_ram.memory[86][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12825_ (.D(_01322_),
    .CLK(net111),
    .Q(\u_cpu.rf_ram.memory[86][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12826_ (.D(_01323_),
    .CLK(net118),
    .Q(\u_cpu.rf_ram.memory[86][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12827_ (.D(_01324_),
    .CLK(net107),
    .Q(\u_cpu.rf_ram.memory[86][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12828_ (.D(_01325_),
    .CLK(net125),
    .Q(\u_cpu.rf_ram.memory[111][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12829_ (.D(_01326_),
    .CLK(net132),
    .Q(\u_cpu.rf_ram.memory[111][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12830_ (.D(_01327_),
    .CLK(net132),
    .Q(\u_cpu.rf_ram.memory[111][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12831_ (.D(_01328_),
    .CLK(net132),
    .Q(\u_cpu.rf_ram.memory[111][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12832_ (.D(_01329_),
    .CLK(net133),
    .Q(\u_cpu.rf_ram.memory[111][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12833_ (.D(_01330_),
    .CLK(net133),
    .Q(\u_cpu.rf_ram.memory[111][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12834_ (.D(_01331_),
    .CLK(net138),
    .Q(\u_cpu.rf_ram.memory[111][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12835_ (.D(_01332_),
    .CLK(net129),
    .Q(\u_cpu.rf_ram.memory[111][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12836_ (.D(_01333_),
    .CLK(net101),
    .Q(\u_cpu.rf_ram.memory[87][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12837_ (.D(_01334_),
    .CLK(net101),
    .Q(\u_cpu.rf_ram.memory[87][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12838_ (.D(_01335_),
    .CLK(net111),
    .Q(\u_cpu.rf_ram.memory[87][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12839_ (.D(_01336_),
    .CLK(net118),
    .Q(\u_cpu.rf_ram.memory[87][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12840_ (.D(_01337_),
    .CLK(net113),
    .Q(\u_cpu.rf_ram.memory[87][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12841_ (.D(_01338_),
    .CLK(net114),
    .Q(\u_cpu.rf_ram.memory[87][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12842_ (.D(_01339_),
    .CLK(net118),
    .Q(\u_cpu.rf_ram.memory[87][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12843_ (.D(_01340_),
    .CLK(net107),
    .Q(\u_cpu.rf_ram.memory[87][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12844_ (.D(_01341_),
    .CLK(net435),
    .Q(\u_cpu.rf_ram.memory[88][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12845_ (.D(_01342_),
    .CLK(net435),
    .Q(\u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12846_ (.D(_01343_),
    .CLK(net436),
    .Q(\u_cpu.rf_ram.memory[88][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12847_ (.D(_01344_),
    .CLK(net437),
    .Q(\u_cpu.rf_ram.memory[88][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12848_ (.D(_01345_),
    .CLK(net435),
    .Q(\u_cpu.rf_ram.memory[88][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12849_ (.D(_01346_),
    .CLK(net436),
    .Q(\u_cpu.rf_ram.memory[88][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12850_ (.D(_01347_),
    .CLK(net436),
    .Q(\u_cpu.rf_ram.memory[88][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12851_ (.D(_01348_),
    .CLK(net435),
    .Q(\u_cpu.rf_ram.memory[88][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12852_ (.D(_01349_),
    .CLK(net334),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12853_ (.D(_01350_),
    .CLK(net286),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12854_ (.D(_01351_),
    .CLK(net286),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12855_ (.D(_01352_),
    .CLK(net286),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12856_ (.D(_01353_),
    .CLK(net334),
    .Q(\u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12857_ (.D(_01354_),
    .CLK(net334),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12858_ (.D(_01355_),
    .CLK(net317),
    .Q(\u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12859_ (.D(_01356_),
    .CLK(net335),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12860_ (.D(_01357_),
    .CLK(net241),
    .Q(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12861_ (.D(_01358_),
    .CLK(net317),
    .Q(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12862_ (.D(_01359_),
    .CLK(net496),
    .Q(\u_cpu.rf_ram.memory[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12863_ (.D(_01360_),
    .CLK(net498),
    .Q(\u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12864_ (.D(_01361_),
    .CLK(net500),
    .Q(\u_cpu.rf_ram.memory[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12865_ (.D(_01362_),
    .CLK(net501),
    .Q(\u_cpu.rf_ram.memory[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12866_ (.D(_01363_),
    .CLK(net501),
    .Q(\u_cpu.rf_ram.memory[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12867_ (.D(_01364_),
    .CLK(net500),
    .Q(\u_cpu.rf_ram.memory[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12868_ (.D(_01365_),
    .CLK(net501),
    .Q(\u_cpu.rf_ram.memory[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12869_ (.D(_01366_),
    .CLK(net496),
    .Q(\u_cpu.rf_ram.memory[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12870_ (.D(_01367_),
    .CLK(net496),
    .Q(\u_cpu.rf_ram.memory[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12871_ (.D(_01368_),
    .CLK(net498),
    .Q(\u_cpu.rf_ram.memory[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12872_ (.D(_01369_),
    .CLK(net500),
    .Q(\u_cpu.rf_ram.memory[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12873_ (.D(_01370_),
    .CLK(net501),
    .Q(\u_cpu.rf_ram.memory[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12874_ (.D(_01371_),
    .CLK(net502),
    .Q(\u_cpu.rf_ram.memory[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12875_ (.D(_01372_),
    .CLK(net500),
    .Q(\u_cpu.rf_ram.memory[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12876_ (.D(_01373_),
    .CLK(net500),
    .Q(\u_cpu.rf_ram.memory[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12877_ (.D(_01374_),
    .CLK(net496),
    .Q(\u_cpu.rf_ram.memory[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12878_ (.D(_01375_),
    .CLK(net496),
    .Q(\u_cpu.rf_ram.memory[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12879_ (.D(_01376_),
    .CLK(net499),
    .Q(\u_cpu.rf_ram.memory[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12880_ (.D(_01377_),
    .CLK(net505),
    .Q(\u_cpu.rf_ram.memory[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12881_ (.D(_01378_),
    .CLK(net507),
    .Q(\u_cpu.rf_ram.memory[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12882_ (.D(_01379_),
    .CLK(net502),
    .Q(\u_cpu.rf_ram.memory[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12883_ (.D(_01380_),
    .CLK(net505),
    .Q(\u_cpu.rf_ram.memory[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12884_ (.D(_01381_),
    .CLK(net505),
    .Q(\u_cpu.rf_ram.memory[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12885_ (.D(_01382_),
    .CLK(net497),
    .Q(\u_cpu.rf_ram.memory[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12886_ (.D(_01383_),
    .CLK(net497),
    .Q(\u_cpu.rf_ram.memory[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12887_ (.D(_01384_),
    .CLK(net499),
    .Q(\u_cpu.rf_ram.memory[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12888_ (.D(_01385_),
    .CLK(net506),
    .Q(\u_cpu.rf_ram.memory[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12889_ (.D(_01386_),
    .CLK(net507),
    .Q(\u_cpu.rf_ram.memory[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12890_ (.D(_01387_),
    .CLK(net507),
    .Q(\u_cpu.rf_ram.memory[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12891_ (.D(_01388_),
    .CLK(net505),
    .Q(\u_cpu.rf_ram.memory[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12892_ (.D(_01389_),
    .CLK(net505),
    .Q(\u_cpu.rf_ram.memory[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12893_ (.D(_01390_),
    .CLK(net497),
    .Q(\u_cpu.rf_ram.memory[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12894_ (.D(_01391_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12895_ (.D(_01392_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12896_ (.D(_01393_),
    .CLK(net438),
    .Q(\u_cpu.rf_ram.memory[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12897_ (.D(_01394_),
    .CLK(net438),
    .Q(\u_cpu.rf_ram.memory[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12898_ (.D(_01395_),
    .CLK(net438),
    .Q(\u_cpu.rf_ram.memory[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12899_ (.D(_01396_),
    .CLK(net437),
    .Q(\u_cpu.rf_ram.memory[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12900_ (.D(_01397_),
    .CLK(net437),
    .Q(\u_cpu.rf_ram.memory[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12901_ (.D(_01398_),
    .CLK(net437),
    .Q(\u_cpu.rf_ram.memory[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12902_ (.D(_01399_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[98][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12903_ (.D(_01400_),
    .CLK(net200),
    .Q(\u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12904_ (.D(_01401_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[98][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12905_ (.D(_01402_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[98][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12906_ (.D(_01403_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[98][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12907_ (.D(_01404_),
    .CLK(net200),
    .Q(\u_cpu.rf_ram.memory[98][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12908_ (.D(_01405_),
    .CLK(net200),
    .Q(\u_cpu.rf_ram.memory[98][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12909_ (.D(_01406_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[98][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12910_ (.D(_01407_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[100][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12911_ (.D(_01408_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[100][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12912_ (.D(_01409_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[100][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12913_ (.D(_01410_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[100][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12914_ (.D(_01411_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[100][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12915_ (.D(_01412_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[100][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12916_ (.D(_01413_),
    .CLK(net176),
    .Q(\u_cpu.rf_ram.memory[100][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12917_ (.D(_01414_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[100][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12918_ (.D(_01415_),
    .CLK(net382),
    .Q(\u_cpu.rf_ram.memory[89][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12919_ (.D(_01416_),
    .CLK(net382),
    .Q(\u_cpu.rf_ram.memory[89][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12920_ (.D(_01417_),
    .CLK(net382),
    .Q(\u_cpu.rf_ram.memory[89][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12921_ (.D(_01418_),
    .CLK(net382),
    .Q(\u_cpu.rf_ram.memory[89][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12922_ (.D(_01419_),
    .CLK(net383),
    .Q(\u_cpu.rf_ram.memory[89][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12923_ (.D(_01420_),
    .CLK(net383),
    .Q(\u_cpu.rf_ram.memory[89][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12924_ (.D(_01421_),
    .CLK(net383),
    .Q(\u_cpu.rf_ram.memory[89][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12925_ (.D(_01422_),
    .CLK(net384),
    .Q(\u_cpu.rf_ram.memory[89][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12926_ (.D(_00025_),
    .CLK(net292),
    .Q(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12927_ (.D(_01423_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12928_ (.D(_01424_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12929_ (.D(_01425_),
    .CLK(net378),
    .Q(\u_cpu.rf_ram.memory[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12930_ (.D(_01426_),
    .CLK(net378),
    .Q(\u_cpu.rf_ram.memory[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12931_ (.D(_01427_),
    .CLK(net378),
    .Q(\u_cpu.rf_ram.memory[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12932_ (.D(_01428_),
    .CLK(net378),
    .Q(\u_cpu.rf_ram.memory[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12933_ (.D(_01429_),
    .CLK(net379),
    .Q(\u_cpu.rf_ram.memory[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12934_ (.D(_01430_),
    .CLK(net378),
    .Q(\u_cpu.rf_ram.memory[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12935_ (.D(_01431_),
    .CLK(net314),
    .Q(\u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12936_ (.D(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(net340),
    .Q(\u_cpu.rf_ram_if.wdata0_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12937_ (.D(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(net340),
    .Q(\u_cpu.rf_ram_if.wdata0_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12938_ (.D(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(net339),
    .Q(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12939_ (.D(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(net339),
    .Q(\u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12940_ (.D(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(net336),
    .Q(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12941_ (.D(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(net336),
    .Q(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12942_ (.D(\u_cpu.cpu.o_wdata0 ),
    .CLK(net336),
    .Q(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12943_ (.D(\u_cpu.rf_ram_if.wtrig0 ),
    .CLK(net285),
    .Q(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12944_ (.D(_01432_),
    .CLK(net281),
    .Q(\u_cpu.rf_ram_if.rdata1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12945_ (.D(_01433_),
    .CLK(net279),
    .Q(\u_cpu.rf_ram_if.rdata0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12946_ (.D(_01434_),
    .CLK(net320),
    .Q(\u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12947_ (.D(\u_cpu.rf_ram_if.rtrig0 ),
    .CLK(net285),
    .Q(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12948_ (.D(_01435_),
    .CLK(net334),
    .Q(\u_cpu.rf_ram_if.rcnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12949_ (.D(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(net341),
    .Q(\u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12950_ (.D(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .CLK(net341),
    .Q(\u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12951_ (.D(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .CLK(net341),
    .Q(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12952_ (.D(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .CLK(net341),
    .Q(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12953_ (.D(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .CLK(net335),
    .Q(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12954_ (.D(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .CLK(net335),
    .Q(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12955_ (.D(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .CLK(net335),
    .Q(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12956_ (.D(\u_cpu.cpu.o_wdata1 ),
    .CLK(net334),
    .Q(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12957_ (.D(\u_cpu.cpu.o_wen0 ),
    .CLK(net279),
    .Q(\u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12958_ (.D(\u_cpu.cpu.o_wen1 ),
    .CLK(net280),
    .Q(\u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _12959_ (.D(\u_scanchain_local.module_data_in[69] ),
    .CLKN(net534),
    .Q(\u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12960_ (.D(_00026_),
    .CLK(net529),
    .Q(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12961_ (.D(_00037_),
    .CLK(net529),
    .Q(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12962_ (.D(_00048_),
    .CLK(net521),
    .Q(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12963_ (.D(_00059_),
    .CLK(net522),
    .Q(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12964_ (.D(_00070_),
    .CLK(net522),
    .Q(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12965_ (.D(_00081_),
    .CLK(net522),
    .Q(\u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12966_ (.D(_00092_),
    .CLK(net519),
    .Q(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12967_ (.D(_00093_),
    .CLK(net519),
    .Q(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12968_ (.D(_00094_),
    .CLK(net520),
    .Q(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12969_ (.D(_00095_),
    .CLK(net520),
    .Q(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12970_ (.D(_00027_),
    .CLK(net517),
    .Q(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12971_ (.D(_00028_),
    .CLK(net517),
    .Q(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12972_ (.D(_00029_),
    .CLK(net517),
    .Q(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12973_ (.D(_00030_),
    .CLK(net516),
    .Q(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12974_ (.D(_00031_),
    .CLK(net518),
    .Q(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12975_ (.D(_00032_),
    .CLK(net515),
    .Q(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12976_ (.D(_00033_),
    .CLK(net514),
    .Q(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12977_ (.D(_00034_),
    .CLK(net516),
    .Q(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12978_ (.D(_00035_),
    .CLK(net514),
    .Q(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12979_ (.D(_00036_),
    .CLK(net514),
    .Q(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12980_ (.D(_00038_),
    .CLK(net513),
    .Q(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12981_ (.D(_00039_),
    .CLK(net513),
    .Q(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12982_ (.D(_00040_),
    .CLK(net513),
    .Q(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12983_ (.D(_00041_),
    .CLK(net513),
    .Q(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12984_ (.D(_00042_),
    .CLK(net513),
    .Q(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12985_ (.D(_00043_),
    .CLK(net516),
    .Q(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12986_ (.D(_00044_),
    .CLK(net516),
    .Q(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12987_ (.D(_00045_),
    .CLK(net516),
    .Q(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12988_ (.D(_00046_),
    .CLK(net517),
    .Q(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12989_ (.D(_00047_),
    .CLK(net519),
    .Q(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12990_ (.D(_00049_),
    .CLK(net519),
    .Q(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12991_ (.D(_00050_),
    .CLK(net519),
    .Q(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12992_ (.D(_00051_),
    .CLK(net521),
    .Q(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12993_ (.D(_00052_),
    .CLK(net521),
    .Q(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12994_ (.D(_00053_),
    .CLK(net521),
    .Q(\u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12995_ (.D(_00054_),
    .CLK(net521),
    .Q(\u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12996_ (.D(_00055_),
    .CLK(net525),
    .Q(\u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12997_ (.D(_00056_),
    .CLK(net525),
    .Q(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12998_ (.D(_00057_),
    .CLK(net525),
    .Q(\u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12999_ (.D(_00058_),
    .CLK(net526),
    .Q(\u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13000_ (.D(_00060_),
    .CLK(net526),
    .Q(\u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13001_ (.D(_00061_),
    .CLK(net525),
    .Q(\u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13002_ (.D(_00062_),
    .CLK(net525),
    .Q(\u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13003_ (.D(_00063_),
    .CLK(net527),
    .Q(\u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13004_ (.D(_00064_),
    .CLK(net527),
    .Q(\u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13005_ (.D(_00065_),
    .CLK(net527),
    .Q(\u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13006_ (.D(_00066_),
    .CLK(net528),
    .Q(\u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13007_ (.D(_00067_),
    .CLK(net528),
    .Q(\u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13008_ (.D(_00068_),
    .CLK(net530),
    .Q(\u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13009_ (.D(_00069_),
    .CLK(net530),
    .Q(\u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13010_ (.D(_00071_),
    .CLK(net530),
    .Q(\u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13011_ (.D(_00072_),
    .CLK(net531),
    .Q(\u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13012_ (.D(_00073_),
    .CLK(net530),
    .Q(\u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13013_ (.D(_00074_),
    .CLK(net530),
    .Q(\u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13014_ (.D(_00075_),
    .CLK(net531),
    .Q(\u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13015_ (.D(_00076_),
    .CLK(net532),
    .Q(\u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13016_ (.D(_00077_),
    .CLK(net532),
    .Q(\u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13017_ (.D(_00078_),
    .CLK(net532),
    .Q(\u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13018_ (.D(_00079_),
    .CLK(net533),
    .Q(\u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13019_ (.D(_00080_),
    .CLK(net533),
    .Q(\u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13020_ (.D(_00082_),
    .CLK(net534),
    .Q(\u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13021_ (.D(_00083_),
    .CLK(net534),
    .Q(\u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13022_ (.D(_00084_),
    .CLK(net534),
    .Q(\u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13023_ (.D(_00085_),
    .CLK(net535),
    .Q(\u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13024_ (.D(_00086_),
    .CLK(net535),
    .Q(\u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13025_ (.D(_00087_),
    .CLK(net535),
    .Q(\u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13026_ (.D(_00088_),
    .CLK(net535),
    .Q(\u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13027_ (.D(_00089_),
    .CLK(net529),
    .Q(\u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13028_ (.D(_00090_),
    .CLK(net537),
    .Q(\u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13029_ (.D(_00091_),
    .CLK(net534),
    .Q(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_2_540 (.ZN(net540));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_2_541 (.ZN(net541));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_2_542 (.ZN(net542));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_2_543 (.ZN(net543));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_2_544 (.ZN(net544));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_2_545 (.ZN(net545));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_2_546 (.ZN(net546));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11995__D (.I(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13038_ (.I(net536),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13039_ (.I(\u_scanchain_local.data_out ),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input4 (.I(io_in[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_in[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout8 (.I(net9),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout9 (.I(net14),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout10 (.I(net14),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout11 (.I(net13),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout12 (.I(net13),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout13 (.I(net14),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout14 (.I(net21),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout15 (.I(net16),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout16 (.I(net20),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout17 (.I(net20),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout18 (.I(net20),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout19 (.I(net20),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout20 (.I(net21),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout21 (.I(net22),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout22 (.I(net42),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout23 (.I(net27),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout24 (.I(net26),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout25 (.I(net26),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout26 (.I(net27),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout27 (.I(net32),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout28 (.I(net30),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout29 (.I(net30),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout30 (.I(net32),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout32 (.I(net41),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout33 (.I(net36),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout34 (.I(net35),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout35 (.I(net36),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout36 (.I(net40),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout38 (.I(net40),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout39 (.I(net40),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout40 (.I(net41),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout41 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net96),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout43 (.I(net44),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(net55),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net46),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout46 (.I(net55),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout47 (.I(net51),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net51),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout49 (.I(net51),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net51),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout51 (.I(net54),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout52 (.I(net54),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net95),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout56 (.I(net60),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net60),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout58 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout59 (.I(net60),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net66),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout61 (.I(net65),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net65),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout63 (.I(net65),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net66),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net76),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout67 (.I(net69),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net69),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout70 (.I(net75),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout71 (.I(net74),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout72 (.I(net74),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout73 (.I(net74),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net76),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(net94),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout77 (.I(net81),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net81),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout79 (.I(net80),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout81 (.I(net83),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout82 (.I(net83),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net93),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout84 (.I(net88),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout85 (.I(net88),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout86 (.I(net88),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net92),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout89 (.I(net92),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout90 (.I(net91),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout91 (.I(net92),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout92 (.I(net93),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net94),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout95 (.I(net96),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout96 (.I(net232),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout97 (.I(net99),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout99 (.I(net104),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout100 (.I(net103),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout101 (.I(net103),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout102 (.I(net103),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout103 (.I(net104),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net110),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout105 (.I(net109),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout106 (.I(net109),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout107 (.I(net109),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout108 (.I(net109),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout109 (.I(net110),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout110 (.I(net123),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout111 (.I(net114),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout112 (.I(net114),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net114),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout114 (.I(net117),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout115 (.I(net117),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout116 (.I(net117),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout117 (.I(net122),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout118 (.I(net120),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout119 (.I(net120),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout120 (.I(net122),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout121 (.I(net122),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout122 (.I(net123),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net142),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout124 (.I(net125),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout125 (.I(net126),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout126 (.I(net130),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout127 (.I(net128),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout128 (.I(net130),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout129 (.I(net130),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout130 (.I(net141),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout131 (.I(net132),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout132 (.I(net135),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout133 (.I(net135),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout134 (.I(net135),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout135 (.I(net140),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout136 (.I(net139),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout137 (.I(net139),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout138 (.I(net140),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout139 (.I(net140),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout140 (.I(net141),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout142 (.I(net162),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout143 (.I(net144),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout144 (.I(net145),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout145 (.I(net150),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout146 (.I(net149),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout147 (.I(net149),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout148 (.I(net150),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout149 (.I(net150),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout150 (.I(net161),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout151 (.I(net158),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout152 (.I(net158),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout153 (.I(net157),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout154 (.I(net157),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout155 (.I(net156),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout156 (.I(net157),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout157 (.I(net158),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout158 (.I(net160),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout159 (.I(net160),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout160 (.I(net161),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout161 (.I(net162),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout162 (.I(net231),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout163 (.I(net169),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout164 (.I(net165),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout165 (.I(net169),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout166 (.I(net168),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout167 (.I(net169),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout168 (.I(net169),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout169 (.I(net180),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout170 (.I(net171),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout171 (.I(net179),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout172 (.I(net178),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout173 (.I(net174),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout174 (.I(net178),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout175 (.I(net176),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout176 (.I(net178),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout177 (.I(net178),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout178 (.I(net179),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout179 (.I(net180),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout180 (.I(net193),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout181 (.I(net184),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout182 (.I(net184),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout183 (.I(net184),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout184 (.I(net185),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout185 (.I(net192),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout186 (.I(net191),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout187 (.I(net188),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout188 (.I(net191),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout189 (.I(net190),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout190 (.I(net191),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout191 (.I(net192),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout192 (.I(net193),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout193 (.I(net230),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout194 (.I(net202),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout195 (.I(net202),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout196 (.I(net201),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout197 (.I(net201),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout198 (.I(net200),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout199 (.I(net200),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout200 (.I(net201),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout201 (.I(net202),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout202 (.I(net206),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout203 (.I(net204),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout204 (.I(net206),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout205 (.I(net206),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout206 (.I(net229),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout207 (.I(net208),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout208 (.I(net211),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout209 (.I(net211),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout210 (.I(net211),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout211 (.I(net216),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout212 (.I(net215),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout213 (.I(net215),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout214 (.I(net215),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout215 (.I(net216),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout216 (.I(net228),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout217 (.I(net219),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout218 (.I(net219),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout219 (.I(net227),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout220 (.I(net221),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout221 (.I(net226),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout222 (.I(net225),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout223 (.I(net225),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout224 (.I(net225),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout225 (.I(net226),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout226 (.I(net227),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout227 (.I(net228),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout228 (.I(net229),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout229 (.I(net230),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout230 (.I(net231),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout231 (.I(net232),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout232 (.I(net512),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout233 (.I(net235),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout234 (.I(net235),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout235 (.I(net245),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout236 (.I(net245),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout237 (.I(net239),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout238 (.I(net239),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout239 (.I(net244),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout240 (.I(net243),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout241 (.I(net243),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout242 (.I(net243),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout243 (.I(net244),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout244 (.I(net245),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout245 (.I(net257),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout246 (.I(net247),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout247 (.I(net251),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout248 (.I(net251),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout249 (.I(net251),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout250 (.I(net251),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout251 (.I(net256),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout252 (.I(net254),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout253 (.I(net254),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout254 (.I(net255),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout255 (.I(net256),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout256 (.I(net257),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout257 (.I(net306),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout258 (.I(net262),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout259 (.I(net262),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout260 (.I(net262),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout261 (.I(net262),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout262 (.I(net267),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout263 (.I(net266),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout264 (.I(net266),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout265 (.I(net266),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout266 (.I(net267),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout267 (.I(net278),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout268 (.I(net272),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout269 (.I(net272),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout270 (.I(net272),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout271 (.I(net272),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout272 (.I(net277),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout273 (.I(net275),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout274 (.I(net275),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout275 (.I(net277),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout276 (.I(net277),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout277 (.I(net278),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout278 (.I(net305),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout279 (.I(net284),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout280 (.I(net284),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout281 (.I(net283),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout282 (.I(net283),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout283 (.I(net284),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout284 (.I(net290),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout285 (.I(net289),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout286 (.I(net289),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout287 (.I(net289),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout288 (.I(net289),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout289 (.I(net290),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout290 (.I(net304),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout291 (.I(net293),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout292 (.I(net293),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout293 (.I(net297),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout294 (.I(net297),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout295 (.I(net297),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout296 (.I(net297),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout297 (.I(net303),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout298 (.I(net302),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout299 (.I(net302),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout300 (.I(net302),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout301 (.I(net302),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout302 (.I(net303),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout303 (.I(net304),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout304 (.I(net305),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout305 (.I(net306),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout306 (.I(net371),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout307 (.I(net312),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout308 (.I(net312),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout309 (.I(net312),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout310 (.I(net311),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout311 (.I(net312),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout312 (.I(net321),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout313 (.I(net314),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout314 (.I(net320),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout315 (.I(net320),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout316 (.I(net318),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout317 (.I(net318),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout318 (.I(net319),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout319 (.I(net320),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout320 (.I(net321),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout321 (.I(net333),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout322 (.I(net326),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout323 (.I(net326),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout324 (.I(net326),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout325 (.I(net326),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout326 (.I(net332),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout327 (.I(net331),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout328 (.I(net331),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout329 (.I(net330),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout330 (.I(net331),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout331 (.I(net332),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout332 (.I(net333),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout333 (.I(net370),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout334 (.I(net338),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout335 (.I(net338),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout336 (.I(net337),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout337 (.I(net338),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout338 (.I(net342),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout339 (.I(net342),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout340 (.I(net341),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout341 (.I(net342),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout342 (.I(net354),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout343 (.I(net347),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout344 (.I(net347),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout345 (.I(net347),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout346 (.I(net347),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout347 (.I(net353),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout348 (.I(net352),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout349 (.I(net352),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout350 (.I(net352),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout351 (.I(net352),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout352 (.I(net353),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout353 (.I(net354),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout354 (.I(net369),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout355 (.I(net357),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout356 (.I(net357),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout357 (.I(net368),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout358 (.I(net363),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout359 (.I(net360),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout360 (.I(net363),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout361 (.I(net363),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout362 (.I(net363),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout363 (.I(net367),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout364 (.I(net366),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout365 (.I(net366),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout366 (.I(net367),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout367 (.I(net368),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout368 (.I(net369),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout369 (.I(net370),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout370 (.I(net371),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout371 (.I(net511),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout372 (.I(net377),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout373 (.I(net377),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout374 (.I(net376),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout375 (.I(net377),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout376 (.I(net377),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout377 (.I(net386),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout378 (.I(net379),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout379 (.I(net385),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout380 (.I(net381),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout381 (.I(net384),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout382 (.I(net384),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout383 (.I(net384),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout384 (.I(net385),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout385 (.I(net386),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout386 (.I(net409),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout387 (.I(net392),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout388 (.I(net392),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout389 (.I(net392),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout390 (.I(net391),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout391 (.I(net392),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout392 (.I(net397),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout393 (.I(net395),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout394 (.I(net395),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout395 (.I(net397),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout396 (.I(net397),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout397 (.I(net408),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout398 (.I(net407),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout399 (.I(net400),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout400 (.I(net407),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout401 (.I(net406),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout402 (.I(net406),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout403 (.I(net405),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout404 (.I(net405),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout405 (.I(net406),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout406 (.I(net407),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout407 (.I(net408),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout408 (.I(net409),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout409 (.I(net451),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout410 (.I(net412),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout411 (.I(net412),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout412 (.I(net418),
    .Z(net412));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout413 (.I(net418),
    .Z(net413));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout414 (.I(net415),
    .Z(net414));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout415 (.I(net417),
    .Z(net415));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout416 (.I(net418),
    .Z(net416));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout417 (.I(net418),
    .Z(net417));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout418 (.I(net428),
    .Z(net418));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout419 (.I(net421),
    .Z(net419));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout420 (.I(net421),
    .Z(net420));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout421 (.I(net427),
    .Z(net421));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout422 (.I(net426),
    .Z(net422));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout423 (.I(net426),
    .Z(net423));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout424 (.I(net426),
    .Z(net424));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout425 (.I(net426),
    .Z(net425));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout426 (.I(net427),
    .Z(net426));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout427 (.I(net428),
    .Z(net427));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout428 (.I(net450),
    .Z(net428));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout429 (.I(net430),
    .Z(net429));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout430 (.I(net434),
    .Z(net430));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout431 (.I(net434),
    .Z(net431));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout432 (.I(net434),
    .Z(net432));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout433 (.I(net434),
    .Z(net433));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout434 (.I(net440),
    .Z(net434));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout435 (.I(net439),
    .Z(net435));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout436 (.I(net439),
    .Z(net436));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout437 (.I(net439),
    .Z(net437));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout438 (.I(net439),
    .Z(net438));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout439 (.I(net440),
    .Z(net439));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout440 (.I(net449),
    .Z(net440));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout441 (.I(net443),
    .Z(net441));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout442 (.I(net443),
    .Z(net442));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout443 (.I(net448),
    .Z(net443));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout444 (.I(net448),
    .Z(net444));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout445 (.I(net447),
    .Z(net445));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout446 (.I(net447),
    .Z(net446));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout447 (.I(net448),
    .Z(net447));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout448 (.I(net449),
    .Z(net448));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout449 (.I(net450),
    .Z(net449));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout450 (.I(net451),
    .Z(net450));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout451 (.I(net510),
    .Z(net451));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout452 (.I(net460),
    .Z(net452));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout453 (.I(net460),
    .Z(net453));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout454 (.I(net455),
    .Z(net454));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout455 (.I(net459),
    .Z(net455));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout456 (.I(net458),
    .Z(net456));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout457 (.I(net458),
    .Z(net457));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout458 (.I(net459),
    .Z(net458));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout459 (.I(net460),
    .Z(net459));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout460 (.I(net470),
    .Z(net460));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout461 (.I(net462),
    .Z(net461));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout462 (.I(net463),
    .Z(net462));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout463 (.I(net469),
    .Z(net463));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout464 (.I(net468),
    .Z(net464));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout465 (.I(net468),
    .Z(net465));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout466 (.I(net467),
    .Z(net466));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout467 (.I(net468),
    .Z(net467));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout468 (.I(net469),
    .Z(net468));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout469 (.I(net470),
    .Z(net469));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout470 (.I(net495),
    .Z(net470));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout471 (.I(net473),
    .Z(net471));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout472 (.I(net476),
    .Z(net472));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout473 (.I(net476),
    .Z(net473));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout474 (.I(net475),
    .Z(net474));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout475 (.I(net476),
    .Z(net475));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout476 (.I(net484),
    .Z(net476));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout477 (.I(net480),
    .Z(net477));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout478 (.I(net480),
    .Z(net478));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout479 (.I(net483),
    .Z(net479));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout480 (.I(net483),
    .Z(net480));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout481 (.I(net483),
    .Z(net481));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout482 (.I(net483),
    .Z(net482));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout483 (.I(net484),
    .Z(net483));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout484 (.I(net494),
    .Z(net484));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout485 (.I(net489),
    .Z(net485));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout486 (.I(net489),
    .Z(net486));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout487 (.I(net489),
    .Z(net487));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout488 (.I(net489),
    .Z(net488));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout489 (.I(net493),
    .Z(net489));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout490 (.I(net492),
    .Z(net490));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout491 (.I(net492),
    .Z(net491));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout492 (.I(net493),
    .Z(net492));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout493 (.I(net494),
    .Z(net493));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout494 (.I(net495),
    .Z(net494));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout495 (.I(net509),
    .Z(net495));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout496 (.I(net498),
    .Z(net496));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout497 (.I(net498),
    .Z(net497));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout498 (.I(net503),
    .Z(net498));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout499 (.I(net503),
    .Z(net499));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout500 (.I(net501),
    .Z(net500));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout501 (.I(net503),
    .Z(net501));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout502 (.I(net503),
    .Z(net502));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout503 (.I(net504),
    .Z(net503));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout504 (.I(net508),
    .Z(net504));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout505 (.I(net506),
    .Z(net505));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout506 (.I(net507),
    .Z(net506));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout507 (.I(net508),
    .Z(net507));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout508 (.I(net509),
    .Z(net508));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout509 (.I(net510),
    .Z(net509));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout510 (.I(net511),
    .Z(net510));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout511 (.I(net512),
    .Z(net511));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout512 (.I(net5),
    .Z(net512));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout513 (.I(net514),
    .Z(net513));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout514 (.I(net515),
    .Z(net514));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout515 (.I(net518),
    .Z(net515));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout516 (.I(net517),
    .Z(net516));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout517 (.I(net518),
    .Z(net517));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout518 (.I(net524),
    .Z(net518));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout519 (.I(net523),
    .Z(net519));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout520 (.I(net523),
    .Z(net520));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout521 (.I(net523),
    .Z(net521));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout522 (.I(net523),
    .Z(net522));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout523 (.I(net524),
    .Z(net523));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout524 (.I(net538),
    .Z(net524));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout525 (.I(net527),
    .Z(net525));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout526 (.I(net527),
    .Z(net526));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout527 (.I(net529),
    .Z(net527));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout528 (.I(net529),
    .Z(net528));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout529 (.I(net537),
    .Z(net529));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout530 (.I(net532),
    .Z(net530));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout531 (.I(net532),
    .Z(net531));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout532 (.I(net536),
    .Z(net532));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout533 (.I(net536),
    .Z(net533));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout534 (.I(net535),
    .Z(net534));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout535 (.I(net536),
    .Z(net535));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout536 (.I(net537),
    .Z(net536));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout537 (.I(net538),
    .Z(net537));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout538 (.I(net1),
    .Z(net538));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_2_539 (.ZN(net539));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11996__D (.I(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11997__D (.I(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__D (.I(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__D (.I(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12000__D (.I(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__D (.I(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__D (.I(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12926__D (.I(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13029__D (.I(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12966__D (.I(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11734__D (.I(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12455__D (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12457__D (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__D (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12659__D (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__I (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__I (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A1 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A2 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__A1 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__I (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__I (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__I (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__I (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__C (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__A2 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__A2 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A3 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__A1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A2 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A2 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A2 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__B (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__A1 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__B (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__B (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A2 (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__A2 (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__A2 (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__A2 (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__A2 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__A1 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__A3 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__B2 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__A3 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__A3 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__B (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__B (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__B (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__I (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__C (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__B2 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__A2 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05816__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__I (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__C (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__C (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__C (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__I (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__I (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__I (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__I (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__B (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__B (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__B (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__I (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__A2 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__I (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__A2 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__A2 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__I (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__I (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__I (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__I (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__I (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__B (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__B (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__B (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__B (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A2 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__A1 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05837__A1 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__A2 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05837__A2 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__I (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__I (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__I (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__I (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__C (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__C (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__C (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__C (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A3 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__A2 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__A2 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__I (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__I (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A4 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__I (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A1 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__I (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__I (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__I (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__I (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05853__I (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05854__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__S0 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__S0 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__S0 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__S0 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__S0 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__S1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__S1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__I (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__I (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__I (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__S1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__S1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__S1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__S1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__S1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__A2 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__I (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__I (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__I (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__I (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__I (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__I (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__I (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__I (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__I (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__I (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__S0 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__S0 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__S0 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__S0 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__S0 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__S0 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__S0 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__I (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__I (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__I (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__I (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__S1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__S1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__S1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__S1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__S1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__A2 (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__B (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__B (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__B (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__B (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__B (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__B (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__B (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__B (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__A2 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__S0 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__S0 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__S0 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__S0 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__S0 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__S1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__S1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__S1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__S1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__S1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A2 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__I (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__I (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05906__I (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__I (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__B (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__B (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__B2 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A1 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__I (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__I (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__I (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__S0 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__S0 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__S0 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__S0 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__S0 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__S1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__S1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__S1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__S1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__S1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__S1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__S1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__S1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__A2 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__S0 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__S0 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__I (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__S0 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__I (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__S0 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__S0 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__S0 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__S0 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__S0 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__S1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__S1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__I (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__S1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__I (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__S1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__S1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__S1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__S1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__S1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__A2 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__I (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__I (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__I (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__I (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__I (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__B (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__B (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__B (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__B (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__B (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__I (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__I (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__I (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__I (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__I (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A1 (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__I (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__S0 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__S0 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__S0 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__S0 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__S0 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__I (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__I (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__I (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__I (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__I (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__S1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__S1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__S1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__S1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__S1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A1 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__A1 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A1 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A1 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A1 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__S0 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__S0 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__S0 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__S0 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__I (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__S0 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__S0 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__S0 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__S0 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__S0 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__S1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__S1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__S1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__S1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__S1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__S1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__S1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__S1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__S1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A2 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__B (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__B (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__B (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__B (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__B (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__I (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__I (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__I (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__I (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__C (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__C (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__I (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__I (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__I (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__C (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__C (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__C (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__C (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__C (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A3 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A1 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A1 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A1 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A1 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__A1 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__I (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__I (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__I (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__I (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__I (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__S0 (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__S0 (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__S0 (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__S0 (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__S0 (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__I (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__I (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__I (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__I (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__I (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__S1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__S1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__S1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__S1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__S1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__A2 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__I (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__I (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__I (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__I (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__I (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__I (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__I (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__I (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__S1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__S1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__S1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__S1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__S1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__A2 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__B (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__B (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__B (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__B (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__B (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__I (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__I (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__I (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__I (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__I (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__S1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__S1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__S1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__S1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__S1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A1 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__A1 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A1 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__A1 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__A1 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__S0 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__S0 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__S0 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__S0 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__S0 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__I (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06189__I (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__I (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__I (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__I (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__S1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__S1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__S1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__S1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__S1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__B (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__B (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__B (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__B (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__B (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__C (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__C (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__C (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__C (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__C (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A2 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__I (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__I (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__I (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__I (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05968__I (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__S0 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__S0 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__S0 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__S0 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__S0 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__I (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__I (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__I (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__I (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__I (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__S1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__S1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__S1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__S1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__S1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__A2 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__A2 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__I (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__I (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__I (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__I (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__I (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05984__A1 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__S0 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__S0 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__S0 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__S0 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__S0 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__S1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__S1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__S1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__S1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__S1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05984__A2 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__A1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06170__A1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__I (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__I (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__I (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__I (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__I (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__S1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__S1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__S1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__S1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__S1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__B (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__B (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__B (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06170__B (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__B (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__B2 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A3 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__S0 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__S0 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__S0 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__S0 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__S0 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__S1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__S1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__S1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__S1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__S1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A1 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A1 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__A1 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__A1 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A1 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__S0 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__S0 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__S0 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__S0 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__S0 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A2 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__A1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__S0 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__S0 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__S0 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__S0 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__S0 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__C (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__C (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__C (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__C (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__C (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A2 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__S0 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__S0 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__S0 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__S0 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__S0 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__S1 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__S1 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__S1 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__S1 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__S1 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A2 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__S0 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__S0 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__S0 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__S0 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__S0 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__S1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__S1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__S1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__S1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__S1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A2 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__B (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__B (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__B (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__B (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__B (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__A2 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__S0 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__S0 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__S0 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__S0 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__S0 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__S1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__S1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__S1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__S1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__S1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__B (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__B (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__B (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__B (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__B (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__C (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__C (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__C (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__C (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__C (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A3 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A1 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A1 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A1 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A1 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A1 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__S0 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__S0 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__S0 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__S0 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__S0 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__S1 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__S1 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__S1 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__S1 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__S1 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A2 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A1 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A1 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A1 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A1 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__A1 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__S0 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__S0 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__S0 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__S0 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__S0 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__S1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__S1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__S1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__S1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__S1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__A2 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__B (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__B (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__B (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__B (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__B (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__S0 (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__S0 (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__S0 (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__S0 (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__S0 (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__A2 (.I(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__S0 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__S0 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__S0 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__S0 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__S0 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__S1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__S1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__S1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__S1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__S1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__A2 (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__B (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__B (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__B (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__B (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__B (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__B2 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__A1 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A1 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A1 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__A1 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__S0 (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__S0 (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__I (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__S0 (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__S0 (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__I (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__S1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__I (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__I (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__S1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__A2 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__S0 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__S0 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__S0 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__S0 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__S0 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__S1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__S1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__S1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__S1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__S1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A2 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__B (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__B (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__B (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__B (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__B (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__S0 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__S0 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__S0 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__S0 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__S0 (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__S1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__S1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__S1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__S1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__S1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__B1 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__S1 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__S1 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__S1 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__S1 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__C (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__C (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__C (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__C (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__C (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A3 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__S0 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__S0 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__S0 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__S0 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__I (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__S0 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__S0 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__S0 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__S1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__S1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__I (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__I (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__I (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__S1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__S1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__S1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__S1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__S1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A2 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A1 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__S0 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__S0 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__S0 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__S1 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__S1 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__S1 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__S1 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__A2 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__B (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__S0 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__S0 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__S0 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__S0 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__S0 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__S1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__S1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__S1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__S1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__S1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__S0 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__S0 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__S0 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__S0 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__S0 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__S1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__S1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__S1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__S1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__S1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__A2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__B (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__S1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__S1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__S1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__S1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__S1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A2 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__A2 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__B2 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__A2 (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__S0 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__S0 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__S0 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__S0 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__S0 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__A2 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A2 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A3 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A2 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A2 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A2 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__S1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__S1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__S1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__S1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__S1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__A2 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__A2 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__B2 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A3 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A2 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__S1 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__S1 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__S1 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__S1 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__S1 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__A2 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__C (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__C (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__C (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__C (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__C (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A2 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__A2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__S1 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__S1 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__S1 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__S1 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__S1 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A2 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__S1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__S1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__S1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__S1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__S1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__A2 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__A2 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A3 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__S1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__S1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__S1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__S1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__S1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A2 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A2 (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__S0 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__S0 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__S0 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__S0 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__S0 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A2 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__B2 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__C (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__C (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__C (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__C (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__C (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__S1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__S1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__S1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__S1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__S1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A2 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A2 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__S0 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__S0 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__S0 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__S0 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__S0 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A2 (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__B1 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A3 (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__S1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__S1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__S1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__S1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__S1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A2 (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A2 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A2 (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A2 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A2 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__S0 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__S0 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__S0 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__S0 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__S0 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A2 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__B2 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A2 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A1 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__S1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__S1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__S1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__S1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__S1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A3 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__A2 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A2 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__A1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__A1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A2 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A2 (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__S1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__S1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__S1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__S1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__S1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__A2 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__B2 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A3 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__S0 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__S0 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__S0 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__S0 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__S0 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__A2 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__A1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__A1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A2 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__S0 (.I(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__S0 (.I(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__S0 (.I(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__S0 (.I(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__S0 (.I(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A2 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A2 (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__A2 (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A3 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__S0 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__S0 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__S0 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__S0 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__S0 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__A2 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A2 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__B2 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A2 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__S1 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__S1 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__S1 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__S1 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__S1 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A2 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__A2 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__A2 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__B2 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A3 (.I(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A2 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__A1 (.I(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A2 (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__S0 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__S0 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__S0 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__S0 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__S0 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A2 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A2 (.I(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__B (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A2 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A2 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__B (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__B (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__B (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__B (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__B (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A2 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__S1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__S1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__S1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__S1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__S1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A2 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A2 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__B2 (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A1 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A2 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__S0 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__S0 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__S0 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__S0 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__S0 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__A2 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A3 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A2 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__S1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__S1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__S1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__S1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__S1 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__A2 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__S0 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__S0 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__S0 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__S0 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__S0 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__S1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__S1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__S1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__S1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__S1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A2 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__A2 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__S1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__S1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__S1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__S1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__S1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A2 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__B1 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A2 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__B2 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__A3 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A2 (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__S0 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__S0 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__S0 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__S0 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__S0 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A1 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A1 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A1 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A1 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A1 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A2 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__B (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__B (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__B (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__B (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__B (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A2 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__A2 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A2 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__S0 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__S0 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__S0 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__S0 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__S0 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A2 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__B1 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__S0 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__S0 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__S0 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__S0 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__S0 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__A2 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A3 (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__S0 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__S0 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__S0 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__S0 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__S0 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A2 (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A2 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__S1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__S1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__S1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__S1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__S1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A2 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A2 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A2 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__B2 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A3 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__S0 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__S0 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__S0 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__S0 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__S0 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A2 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__S1 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__S1 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__S1 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__S1 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__S1 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__A2 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A2 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06467__A2 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A2 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A2 (.I(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A2 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A2 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A1 (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A2 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A2 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__A3 (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A2 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A2 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A2 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A2 (.I(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__B1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A2 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__B2 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A3 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A2 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A2 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A2 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__A2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A2 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A2 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A3 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A2 (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A2 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A2 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__A2 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06533__A2 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A2 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A2 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__B2 (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__A3 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A2 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A2 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A2 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A2 (.I(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__B (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A2 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A1 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A2 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A2 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A2 (.I(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__A1 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06567__A2 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A3 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A2 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A2 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__B1 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A2 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__A2 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__B1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__B2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A3 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A2 (.I(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A2 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A2 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A2 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A3 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__A2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A2 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A2 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A2 (.I(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A2 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A2 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A3 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A2 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A2 (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A2 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A2 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__B (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__A2 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__A2 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__B2 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A2 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A3 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A2 (.I(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__A2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A2 (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A2 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06675__A2 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__B1 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__B2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A3 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__A2 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A2 (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__A2 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__A2 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__A3 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A2 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__A2 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__A2 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A2 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A2 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A3 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A2 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A2 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A2 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__B (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A1 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A2 (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A2 (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A2 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A3 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A2 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A2 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A2 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A2 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__B1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__B2 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A3 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A2 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__B1 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A2 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A2 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A2 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A3 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__A2 (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A2 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__A2 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A2 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A3 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A2 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__A2 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__I (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__B (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__I (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A2 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__B1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__B (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__B (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__B2 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__A2 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A1 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A2 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__A3 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__I1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__B2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__A2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A1 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A1 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A1 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__C (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A1 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A1 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A1 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__I (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__A1 (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__B (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A2 (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__B (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__A1 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A1 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A3 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A4 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A4 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A2 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A2 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A2 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__C (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__B2 (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A2 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__A1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A2 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A2 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__B2 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A2 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A2 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__A1 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__I (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__B (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__B (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__I (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__I (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A2 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__A1 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__A1 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A2 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__I (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__I (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A2 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A2 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__A1 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A2 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A2 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A2 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A2 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A2 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A2 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__B1 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__C (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A2 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A2 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A1 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__A1 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__A1 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__A1 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__B1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A2 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__I (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A2 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A2 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__A1 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__B2 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06915__A2 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__C (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__I1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A3 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__C (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__B (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__I (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__A1 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A1 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__C (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A3 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A2 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__I0 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__B (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A2 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__I1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__I (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__A2 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A2 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A2 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A2 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A2 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A2 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A2 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A2 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A2 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A1 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A1 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A1 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__I (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A3 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__C (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A1 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__C (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__A2 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A1 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__B (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__I (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__A2 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__I (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A2 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__I (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__I (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A2 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A2 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__B1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__B1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__C1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__B (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__I (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__I (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__I (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__I (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__B (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A2 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__C (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__B (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A2 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__A2 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A2 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A2 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A2 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A3 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__A1 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A1 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__I1 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__S (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__S (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__S (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__S (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__S (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A1 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__I (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__I (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__I (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__I (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__S (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__S (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__S (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__S (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__S (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__S (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__S (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__S (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__S (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__S (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__S (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__S (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__S (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__S (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__S (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A1 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A1 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__S (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__S (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__S (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A1 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A1 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A1 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A1 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A1 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A2 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A2 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__B2 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A2 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A3 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A2 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A2 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__A2 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__I (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A1 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A1 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__C (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__B (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__I (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__I (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__B1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__A1 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__A1 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A1 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__S (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__S (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A1 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A1 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__I (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__I (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__I (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A1 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__I (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__S (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__S (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__I (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A1 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__B (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__B (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__B (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__I (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A1 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A1 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__A1 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__A1 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__A1 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A1 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__S (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A1 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A1 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A1 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__B1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__B1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__B1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__B1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__B1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__S (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__S (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__A4 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07156__A3 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__I (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__I (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__I (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__B1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__B1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__B1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__B1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__B1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A1 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A1 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A1 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A1 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A3 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__I (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__B2 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A3 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A3 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A2 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A2 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A3 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__C (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__B (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__C (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__B1 (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__B1 (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__B1 (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__B1 (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__B1 (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__B2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A4 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A2 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A2 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__B (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__B (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__B (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__B1 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__B1 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__B1 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__B1 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__B1 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A1 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A1 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A1 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A1 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A4 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__C (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A3 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A4 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A1 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__B (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__I (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A2 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__B (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__B (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A1 (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__A2 (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A1 (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__B (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__B (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A1 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A1 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A1 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__A1 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A3 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__A3 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A2 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__B (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A3 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__B (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__C (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__I (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A2 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__I (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__B1 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A1 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A1 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A1 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A1 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__S (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__I (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A2 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A2 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__I (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A1 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A2 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A2 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__A1 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A2 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__A1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__A1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A1 (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__I (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__I (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__I (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__A1 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A1 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A1 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__A1 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__A1 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A1 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A1 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__A1 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A1 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A1 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__A1 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__A1 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A2 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__A2 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__I (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__I (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__I (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__I (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__I (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__I (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__I (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__I (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__I (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__I (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__I (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__I (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__I (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__I (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A1 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A1 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A1 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A1 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__A2 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A2 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__A2 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__I (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__I (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__I (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__I (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__I (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__I (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__I (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__I (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__I (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__I (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__I (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__I (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__I (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__I (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__I (.I(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__I (.I(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__I (.I(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__I (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__I (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__I (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__I (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__I (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__I (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__I (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__I (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__I (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__I (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A2 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__A2 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__A2 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A2 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A2 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__A2 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__I (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__I (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__I (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__I (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__I (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__I (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__I (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__I (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__I (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__I (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__I (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__I (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__I (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__I (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A1 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A1 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A1 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A1 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__A2 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__I (.I(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__I (.I(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__I (.I(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__I (.I(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__I (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__I (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__I (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__I (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__I (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__I (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__I (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__I (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__I (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__I (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__I (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__I (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__I (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__I (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__I (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__I (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__I (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__I (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__I (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__I (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__I (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__I (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__I (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A1 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__A1 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A1 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__I (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__I (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__I (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__I (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__I (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__I (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__I (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__I (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__I (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__I (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__I (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__I (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__I (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__I (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A2 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A2 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A2 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__I (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A2 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A2 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A3 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A3 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A2 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A4 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__I (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__I (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__I (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A2 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A2 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A1 (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A1 (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A1 (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A1 (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A1 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A1 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A1 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__I (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A1 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A1 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A1 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A2 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A2 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A2 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A2 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A2 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A2 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A2 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A2 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A2 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A2 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__A1 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A1 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A1 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A1 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__I (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A1 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A1 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A1 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A2 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A2 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A2 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A2 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A1 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A1 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A1 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__A1 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A1 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__A1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A2 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__I (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__I (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__I (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A2 (.I(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__I (.I(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__I (.I(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__I (.I(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A2 (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A2 (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A2 (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A2 (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__A2 (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A1 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A1 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__I (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__A2 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A2 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A1 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A1 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A2 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A2 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A2 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A2 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A2 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A2 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__I (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__A2 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A2 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__A2 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A2 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A2 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A2 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A2 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__I (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A2 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A2 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A2 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A3 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A3 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A4 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A4 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A4 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A1 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A2 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A2 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A2 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A2 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A2 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A2 (.I(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A2 (.I(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A2 (.I(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__A2 (.I(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__A2 (.I(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A1 (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A1 (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A1 (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__I (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A1 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__I (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__I (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__I (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__A2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__A2 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A2 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A2 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A2 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A2 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A2 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A2 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A2 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__A2 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__A2 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A1 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A1 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A1 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A1 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A1 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A2 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__A1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__I (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A2 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A2 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A2 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A2 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A2 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A2 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A2 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A2 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A2 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A1 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A2 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A2 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__A2 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__A2 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A2 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A1 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A1 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A1 (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A1 (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A1 (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__I (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A1 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A1 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A1 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__I (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A1 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__I (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__I (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__I (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A2 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__I (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A2 (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A2 (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A2 (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A2 (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A2 (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A1 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A1 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__I (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__A2 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A2 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A2 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A2 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A2 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A1 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A1 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A1 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A1 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A1 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A2 (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__I (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__I (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__I (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__A2 (.I(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A2 (.I(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A2 (.I(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__A2 (.I(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A2 (.I(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A1 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A1 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A1 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A1 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A1 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A1 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A1 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A1 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A1 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A1 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A1 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A1 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A1 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A1 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A2 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A1 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A1 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__I (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A2 (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__I (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__I (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__I (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A1 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__A1 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A1 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A2 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A2 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A2 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__B (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__I (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__I (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__I (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__I (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__I (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__B (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__A1 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A1 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A1 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__B (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A1 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A1 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A2 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A2 (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__C (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A2 (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A2 (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__B2 (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A3 (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A1 (.I(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__I (.I(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__B (.I(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__A1 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__A2 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A2 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A2 (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__I (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__I (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__I (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A2 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A2 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__I (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__I (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__I (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__I (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__I (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A1 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A1 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A1 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A2 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__I (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__I (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__I (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__I (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__I (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__I (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__I (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__I (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__I (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__I (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__I (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A1 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A1 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A1 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A1 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A1 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__I (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__I (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__I (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__I (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__I (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A1 (.I(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A1 (.I(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A1 (.I(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A1 (.I(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A1 (.I(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__I (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__I (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__I (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__I (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A1 (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__A1 (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A1 (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__I (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__I (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__I (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__I (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__I (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__I (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__I (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__I (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__I (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__I (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__I (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__I (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__I (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__I (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__I (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__I (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__I (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__I (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A2 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A2 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__I (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A1 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__I (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__I (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A2 (.I(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A2 (.I(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A2 (.I(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A2 (.I(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A2 (.I(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A2 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A2 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A2 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A2 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A2 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A2 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A2 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A2 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A2 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A1 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A1 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A2 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A2 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A2 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A2 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A2 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A2 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__I (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__I (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__I (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A2 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A2 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A2 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A2 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A1 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A1 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A1 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A1 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A1 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A1 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A1 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A1 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A1 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__A1 (.I(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A1 (.I(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A1 (.I(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A1 (.I(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A1 (.I(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__I (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__I (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__I (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A2 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A2 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A2 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A2 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A2 (.I(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A2 (.I(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A2 (.I(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A2 (.I(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A2 (.I(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A1 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A2 (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__I (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__I (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__I (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A2 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A2 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A2 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A2 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A2 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A2 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__A2 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A2 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A2 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A2 (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A1 (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A2 (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A2 (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__I (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A2 (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__I (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__I (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__I (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A2 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A2 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A2 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A2 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A2 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A2 (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__I (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__I (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__I (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A2 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A2 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A2 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A2 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A2 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A2 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A2 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A2 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A2 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A2 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A2 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A2 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A2 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A2 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A2 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A2 (.I(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__I (.I(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__I (.I(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__I (.I(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A2 (.I(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A2 (.I(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A2 (.I(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A2 (.I(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A2 (.I(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__A2 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A2 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A2 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A2 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A2 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A2 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A2 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A2 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__A2 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A2 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A1 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A1 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A1 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A1 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__A1 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A2 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__I (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__I (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__I (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A2 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A2 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A2 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__A2 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__I (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__I (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__I (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A2 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A2 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A2 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A2 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A2 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__I (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__I (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__I (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A2 (.I(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A2 (.I(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A2 (.I(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A2 (.I(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A2 (.I(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A1 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A1 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A1 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A2 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A2 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A2 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A2 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A2 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A2 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A2 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A2 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A2 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A2 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A2 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__A1 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A1 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A1 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A1 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A1 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A2 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__I (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__I (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__I (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A2 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A2 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A2 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A2 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A1 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A1 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A1 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A1 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A1 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A2 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A2 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A2 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__A2 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A2 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A1 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A1 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A1 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A1 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A1 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A1 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__I (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__I (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__I (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A2 (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A2 (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A2 (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A2 (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A2 (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A2 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A2 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A2 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A2 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A2 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A2 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A2 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A2 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__I (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__I (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__I (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A2 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A2 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A2 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A2 (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A2 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A2 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A2 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A2 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A2 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A2 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A2 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A2 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A2 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A2 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__I (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A2 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A2 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A2 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A2 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__A1 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__A1 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__A1 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A1 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__I (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11491__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__I (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__A1 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A1 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A1 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__A1 (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__A1 (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__A1 (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A1 (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__I (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A1 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A1 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__A1 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A1 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__I (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__A1 (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__A1 (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__A1 (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__A1 (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__I (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A1 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A1 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A1 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A1 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A1 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11539__A1 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__A1 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__A1 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__I (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A1 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A1 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A1 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A1 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A1 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__I (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A1 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A1 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A2 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A2 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A2 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A2 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A2 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A2 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A2 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A2 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A2 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__I (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__I (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__I (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A2 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A2 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A2 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A2 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A2 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A2 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A2 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A2 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A2 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__I (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__I (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__I (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__I (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__I (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A1 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A1 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A1 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__A1 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A2 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A2 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A2 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A2 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__A2 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__I (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__I (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__I (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__I (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__I (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__I (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__I (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__I (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__I (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A1 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A1 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A1 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A1 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A1 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__I (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__I (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__I (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__I (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__I (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__I (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__I (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__I (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__I (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__I (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__I (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__I (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__I (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__I (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__I (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__I (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A2 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A2 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A2 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A2 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A2 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A2 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A2 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A2 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A2 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A2 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A2 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A2 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__I (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__I (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__I (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A2 (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A2 (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A2 (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A2 (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A2 (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A2 (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A2 (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A2 (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A2 (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A2 (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__I (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__I (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__I (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__A2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__A2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__A2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__I (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A2 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A1 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A1 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A1 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__I (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__I (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__I (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A2 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A2 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A2 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A2 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A2 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A2 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A1 (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A1 (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A1 (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A1 (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A1 (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A1 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A1 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A1 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A1 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A2 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__I (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__I (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__I (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A2 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__I (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__I (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__I (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A2 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A2 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A2 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A2 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A2 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A2 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A2 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A2 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A2 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A2 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A2 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A2 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A2 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__I (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A1 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A1 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A1 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A1 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A1 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A1 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A1 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A1 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A1 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A1 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A1 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A1 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A2 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__I (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__I (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__I (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A2 (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A2 (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A2 (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A2 (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A2 (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A2 (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__I (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__I (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__I (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__I (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__I (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__I (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A1 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A1 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A1 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A1 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A1 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A1 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A2 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A2 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A2 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A2 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A2 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A2 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A2 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A2 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A2 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A2 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A2 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A2 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__I (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__I (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__I (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A2 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A2 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A2 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A2 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A2 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A2 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__I (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__I (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__I (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A2 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A2 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A2 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A2 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A2 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A2 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A2 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A2 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A2 (.I(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A1 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A1 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A1 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__I (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A2 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A2 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A2 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A2 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A2 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A1 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__A1 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A1 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A1 (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A1 (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A1 (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A1 (.I(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A1 (.I(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A1 (.I(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A1 (.I(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A1 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__A1 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A1 (.I(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__A1 (.I(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__A1 (.I(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A1 (.I(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A1 (.I(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A2 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A2 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A2 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A2 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A2 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A1 (.I(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A1 (.I(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A1 (.I(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A1 (.I(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A1 (.I(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A1 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A1 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A1 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A1 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A1 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A1 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A1 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A1 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A1 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A1 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A1 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A1 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A1 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A2 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A2 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A2 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A2 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A2 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A2 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A2 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A2 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A2 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A2 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__A2 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A2 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__A2 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A2 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__A2 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A2 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__A2 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A2 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A2 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A2 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A2 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A2 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A2 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__I (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__I (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__I (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__I (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__I (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A2 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__I (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__I (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__I (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A1 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A1 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A1 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A1 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__I (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__I (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__I (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__I (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__I (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__I (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__I (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__I (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__I (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__I (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A1 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A1 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A1 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__A1 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A1 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A1 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A1 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A1 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A1 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A2 (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A2 (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A2 (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A2 (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A2 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__I (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__I (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__I (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A2 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A2 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A2 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A2 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A2 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__I (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__I (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__I (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A2 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09328__A2 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A2 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A2 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A2 (.I(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__I (.I(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__I (.I(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__I (.I(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A2 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A2 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A2 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__A2 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A1 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A1 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A2 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A1 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__A1 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__B (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A1 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A1 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__B (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A2 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A1 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A1 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A1 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A2 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A2 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A2 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__A2 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A1 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A1 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A1 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A1 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A2 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A2 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A2 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A2 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A2 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A2 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A2 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A2 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A2 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A2 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A1 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A1 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__A1 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A1 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A1 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A2 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A2 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A2 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A2 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A2 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A2 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__A2 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A2 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A2 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A2 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A2 (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__I (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__I (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__I (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A2 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A2 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A2 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A1 (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A1 (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A1 (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A1 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A1 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A1 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A1 (.I(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A1 (.I(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A1 (.I(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A1 (.I(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__I (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__I (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A2 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A2 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A2 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A2 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A2 (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A2 (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A2 (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A2 (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A2 (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A2 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A2 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A2 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A2 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A2 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__I (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__I (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__I (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A2 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A2 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A2 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A2 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__I (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__I (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__I (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A2 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A2 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A2 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A2 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__I (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__I (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09642__I (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A2 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A2 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A2 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09655__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A2 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__I (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__I (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__I (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A1 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A1 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A1 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A1 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A1 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A1 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A1 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A2 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__I (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__I (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__I (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A2 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A2 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A2 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A2 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A2 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A2 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A2 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A2 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A2 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A2 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A2 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A2 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A2 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A2 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__I (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__A2 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A1 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A2 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A2 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__A2 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A2 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A2 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A2 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__B (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__I (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__I (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__I (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__I (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A2 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A2 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A2 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A2 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__A2 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A2 (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A2 (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__I (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__C (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__I (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__I (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__I (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__I (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__I (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__B1 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__B1 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__B1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A2 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__B1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__B1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__B1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A2 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A2 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__A2 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A2 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__A2 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__B1 (.I(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__B1 (.I(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__B1 (.I(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__B1 (.I(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__B1 (.I(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A2 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A2 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A2 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A2 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A2 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__B1 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A2 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__B1 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A2 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__B (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__A2 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__I (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__I (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__I (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A2 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A2 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A2 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A2 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A2 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__I (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__I (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__I (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__I (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A1 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A1 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__I (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__I (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__C (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__C (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__I (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__S (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__S (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__S (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__I (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A1 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__S (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__S (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__S (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__I (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__S (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A1 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__S (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A1 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A1 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A1 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A4 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__I (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A1 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__B (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__B2 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A2 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A2 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A2 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A1 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__A1 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__B1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__I (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__B1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__B (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__I (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__I (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A1 (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A2 (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__B1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A2 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A2 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A1 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A1 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__B1 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A2 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A2 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__B (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__B (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__B (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__I (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__C (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A1 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A1 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__B1 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__B1 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__I (.I(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__A2 (.I(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__I (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__I (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A1 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A3 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A2 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A2 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__I (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A2 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__B1 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__I (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A1 (.I(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__I (.I(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__A2 (.I(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A2 (.I(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__B (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__I (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A3 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A1 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__I (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A4 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__B1 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__B1 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A2 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A2 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A2 (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__B2 (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A1 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A1 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__I (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A2 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A1 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A1 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__I (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A2 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A1 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A1 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A1 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__A1 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A1 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__I (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A1 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__C (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__B (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__A2 (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__I (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A2 (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__A1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__B2 (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__B2 (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__B2 (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__I (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A2 (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__C2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__B2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A3 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A2 (.I(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A1 (.I(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A1 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__B2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__B (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__A3 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A2 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A3 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A2 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A2 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A3 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A2 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A2 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__A2 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__A2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__B2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A1 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A1 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__A1 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A1 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A2 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A2 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A2 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A2 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__B2 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A1 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__B (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__B (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__C (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__B (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A1 (.I(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A2 (.I(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__C (.I(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__I (.I(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A2 (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A2 (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A2 (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A2 (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A1 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A1 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__B (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__B1 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__B (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__I (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__I (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__I (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A1 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__B (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__C (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__B (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__C2 (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__C2 (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__B2 (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__B2 (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__B (.I(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__B (.I(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A1 (.I(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__C (.I(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A2 (.I(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__B2 (.I(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A2 (.I(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A1 (.I(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A1 (.I(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A1 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A1 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__B2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A2 (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__B2 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A3 (.I(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A1 (.I(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A2 (.I(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A2 (.I(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A2 (.I(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__A2 (.I(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A1 (.I(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__I (.I(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A2 (.I(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__C (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__I (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__B (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__B (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A3 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__C (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A2 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A2 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__B2 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__C (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__I (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__C (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__C (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A1 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__I (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__B1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__B (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__B1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__B (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__B2 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A1 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A1 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A1 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A1 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A1 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A1 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A2 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A2 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A2 (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A2 (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__I (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__B (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__B (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__B (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__I (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__C (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A2 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A2 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__B (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__I (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A2 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A1 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__B2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__I (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A2 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A2 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A1 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A2 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A2 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A1 (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__A1 (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__B2 (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__C (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__B (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A1 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__C (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__B (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A2 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__I (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__A1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A2 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__B2 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__B1 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A1 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A2 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A1 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A1 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A2 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A2 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A1 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__I (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A1 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A3 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A2 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__A2 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__C1 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__B1 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A2 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__B2 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A1 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A1 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A2 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__B2 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A2 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__B1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__B1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__I (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A2 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__B1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__C (.I(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A1 (.I(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__C (.I(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A2 (.I(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__B2 (.I(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A2 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__B2 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__B (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__B (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__B (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__B (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__C (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__I (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A1 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A2 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A1 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__B1 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A1 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A2 (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A2 (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__C (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A4 (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__B (.I(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__B2 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__B2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__B (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A2 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A2 (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__B2 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__B (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A2 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A1 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A1 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__I (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__A1 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__B1 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__A4 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A3 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A2 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A1 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A3 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A1 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A1 (.I(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__B (.I(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A1 (.I(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A3 (.I(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__B (.I(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__B2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A1 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__B (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__B1 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__C2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__C2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__A1 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A1 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__S (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__S (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__S (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A2 (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__B1 (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__B1 (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__C1 (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A2 (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__B (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__C (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__A1 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A3 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__B1 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__C (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__C (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A2 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A2 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__B2 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__B (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A2 (.I(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__B2 (.I(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__B (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__C (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__I (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__I (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__C (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A2 (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A3 (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__C (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A1 (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__B (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__B2 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__B (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A1 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__A1 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A1 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A1 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A2 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__I (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__I (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__I (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A2 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A2 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A2 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A2 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A2 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__A1 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A1 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A1 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A1 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A1 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__A1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A1 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A1 (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A1 (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A1 (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A1 (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__A1 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A1 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__A1 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A1 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A2 (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__B2 (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__C (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A3 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A2 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A2 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A2 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__B (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__I (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__A2 (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A2 (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__C (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A1 (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A2 (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__B (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__B (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__B (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__B (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A1 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__I (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A2 (.I(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__B (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A1 (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__B2 (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__C2 (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__B2 (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A2 (.I(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__B (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A2 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A2 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A2 (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__B1 (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__B (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__C (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__C (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A2 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__B (.I(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A2 (.I(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A1 (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A1 (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__B (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A1 (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__A2 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A1 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A1 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A1 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A1 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A2 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__B1 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__B1 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__B2 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__B1 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__C1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__B2 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__A3 (.I(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A2 (.I(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A2 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A3 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__A2 (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A2 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A2 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A2 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A2 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__B (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__B1 (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__B1 (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A3 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A1 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__B2 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__A1 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A1 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A1 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__C1 (.I(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__B1 (.I(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A2 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A2 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A2 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__A1 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__C (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A2 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__B (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__A1 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A1 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A2 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A1 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A2 (.I(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__C1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A2 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__B1 (.I(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A1 (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__B2 (.I(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A1 (.I(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A2 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A2 (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A2 (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__B (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__B (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__I (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__B (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__I (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__B (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__B (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__B (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A1 (.I(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A1 (.I(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__B (.I(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A2 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A2 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A1 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A1 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__B (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__B1 (.I(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__B (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A2 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__C (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A2 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A2 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__C (.I(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A2 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__B2 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A2 (.I(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__C (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A2 (.I(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A3 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__C (.I(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A2 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__I (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__I (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__I (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A2 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A2 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A2 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A2 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A2 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__I (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__S (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__S (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__S (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__S (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__S (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__S (.I(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__S (.I(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__S (.I(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__S (.I(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__S (.I(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__S (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__S (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__S (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__S (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__S (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__S (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__S (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__S (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__S (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__S (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__B (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__I1 (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A2 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A2 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A2 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A2 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__A2 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A2 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A2 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A2 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A2 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__A2 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A2 (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__A2 (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A2 (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__I (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__I (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__A1 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A2 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A2 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A2 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__A2 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__I (.I(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__I (.I(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__I (.I(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__I (.I(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__B1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__B1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__I (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__I (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__I (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__B1 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__B1 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__B1 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__B1 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__B1 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__A2 (.I(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__A2 (.I(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A2 (.I(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__A2 (.I(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A2 (.I(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A2 (.I(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A2 (.I(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A2 (.I(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A2 (.I(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__A2 (.I(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__B1 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__B1 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__B1 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__B1 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__B1 (.I(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__B1 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__B1 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__B1 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__B1 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__B1 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__B1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__B1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__B1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__B1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__B1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__A2 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A2 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A2 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A2 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__B1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__B1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__B1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__B1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__B1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__B2 (.I(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__I (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__I (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__I (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A2 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A2 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A2 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A2 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A2 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A2 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A2 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A2 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A2 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A2 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A2 (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__I (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__I (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__I (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A2 (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A2 (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A2 (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A2 (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A2 (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A1 (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A1 (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A1 (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A1 (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__A2 (.I(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__I (.I(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__I (.I(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__I (.I(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A2 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A2 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__A2 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A2 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A2 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A2 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A2 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A2 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__A2 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A2 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__I (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__I (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__I (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__I (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__I (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__I (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A1 (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__A1 (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A1 (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__A1 (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A2 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A2 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__A2 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__A2 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A2 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__I (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__I (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__I (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__I (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__I (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__I (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__I (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__I (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__I (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__I (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A1 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A1 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A1 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A1 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A1 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11227__I (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__I (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__I (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__I (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__I (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A1 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__A1 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__A1 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A1 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A1 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__I (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__I (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__I (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__I (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__I (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__A1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__A2 (.I(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A2 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__B1 (.I(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A2 (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__B (.I(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A2 (.I(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__B (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__A3 (.I(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__B1 (.I(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__A2 (.I(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__I (.I(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__I (.I(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__I (.I(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A2 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A2 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A2 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A2 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A2 (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A2 (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__I (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__I (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__I (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A2 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A2 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A2 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A2 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A2 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__A2 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A2 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A2 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__A2 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__A2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__A2 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__I (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__I (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__I (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A2 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A2 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__A2 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A2 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A2 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__A2 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__A2 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A2 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A2 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__A2 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A2 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__A2 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__A2 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A2 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A2 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A2 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__I (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__I (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__I (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A2 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A2 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A2 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A2 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A2 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__A2 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__A2 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A2 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A2 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A2 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A1 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A1 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A1 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A1 (.I(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A1 (.I(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A1 (.I(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A1 (.I(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A1 (.I(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A1 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A1 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A1 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A1 (.I(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A1 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A1 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A1 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A1 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A1 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A1 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A1 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A1 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__A1 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__A1 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A1 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A1 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A1 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A1 (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A1 (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A1 (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A1 (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__A1 (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__S (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__S (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__I (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__I (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__I (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__S (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__S (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__S (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__S (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__S (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__S (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__S (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__S (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__S (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__S (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A2 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__I (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__I (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__I (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A2 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A2 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A2 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A2 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A2 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A2 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__I (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__I (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__I (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A2 (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__I (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__I (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__I (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__A2 (.I(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A2 (.I(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A2 (.I(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A2 (.I(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A2 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A1 (.I(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A1 (.I(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A1 (.I(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A1 (.I(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A2 (.I(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__I (.I(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__I (.I(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__I (.I(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__A2 (.I(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__A2 (.I(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A2 (.I(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A2 (.I(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A2 (.I(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A1 (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A1 (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A1 (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A1 (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A1 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A1 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A1 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A1 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A1 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__A2 (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__A2 (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A2 (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A2 (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A2 (.I(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__A1 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A1 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A1 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__A1 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A2 (.I(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__I (.I(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__I (.I(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__I (.I(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__I (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__I (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__I (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__A2 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A2 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A2 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A2 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A2 (.I(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A2 (.I(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A2 (.I(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__A2 (.I(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A2 (.I(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__A2 (.I(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A2 (.I(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A2 (.I(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A2 (.I(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__A2 (.I(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A2 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__I (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__I (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__I (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A2 (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A2 (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A2 (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A2 (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A2 (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A2 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A2 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A2 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A2 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A2 (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__A2 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__I (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__I (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__I (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A2 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__A2 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__A2 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A2 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A2 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A2 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A1 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A1 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A1 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__A1 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A1 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A1 (.I(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A1 (.I(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A1 (.I(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A1 (.I(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A1 (.I(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A1 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__A1 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__A1 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A1 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A1 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A1 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A1 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A1 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A1 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__A1 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A1 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A1 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A1 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A1 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A1 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A1 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A1 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A1 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A1 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A1 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A1 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A1 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A1 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A2 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A2 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A2 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__A2 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A2 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__A2 (.I(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A2 (.I(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__I (.I(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__I (.I(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__I (.I(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A2 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__A2 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A2 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A2 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A2 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A2 (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A2 (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A2 (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__A2 (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A2 (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A2 (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__I (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__I (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__I (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A2 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__I (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__I (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__I (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A2 (.I(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A2 (.I(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A2 (.I(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A2 (.I(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A2 (.I(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A2 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A2 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A2 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A2 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A2 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A2 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A2 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A2 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A2 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A2 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11297__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__A2 (.I(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__I (.I(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__I (.I(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11207__I (.I(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A1 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A1 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A1 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__A1 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__A2 (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A2 (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__A2 (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A2 (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A2 (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A1 (.I(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A1 (.I(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A1 (.I(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A1 (.I(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__A1 (.I(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A1 (.I(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A1 (.I(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A1 (.I(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A1 (.I(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__A1 (.I(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A1 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A1 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A1 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__A1 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A1 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__A1 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A1 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A1 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A1 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A2 (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__I (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__I (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__I (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A2 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A2 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A2 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A2 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A2 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A2 (.I(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__I (.I(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__I (.I(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__I (.I(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A2 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A2 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A2 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A2 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A2 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A2 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__A2 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A2 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A2 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A2 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A2 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__I (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__I (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A2 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A2 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A2 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A2 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11297__A2 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A2 (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A2 (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A2 (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A2 (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A2 (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__A1 (.I(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A1 (.I(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__A1 (.I(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A1 (.I(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A1 (.I(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A2 (.I(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__I (.I(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__I (.I(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__I (.I(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A1 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__A1 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__A1 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A1 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A1 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A1 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A1 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A1 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__A1 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A1 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A1 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11433__A1 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A1 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A1 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__A1 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A1 (.I(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A1 (.I(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A1 (.I(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A1 (.I(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A1 (.I(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A1 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A1 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A1 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__A1 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A1 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A1 (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11439__A1 (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A1 (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A1 (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__A1 (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A1 (.I(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__A1 (.I(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A1 (.I(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A1 (.I(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A1 (.I(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__B (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__S (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__I (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A2 (.I(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__I (.I(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__I (.I(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__I (.I(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A2 (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A2 (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__A2 (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A2 (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A2 (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A2 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A2 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__A2 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__A2 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11390__A2 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A2 (.I(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__I (.I(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__I (.I(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__I (.I(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A2 (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A2 (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A2 (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__A2 (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__A2 (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A2 (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A2 (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A2 (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A2 (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__A2 (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A2 (.I(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A2 (.I(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A2 (.I(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A2 (.I(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A2 (.I(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__A2 (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__I (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__I (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__I (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A2 (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11433__A2 (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A2 (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__A2 (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A2 (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__A2 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11439__A2 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A2 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__A2 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__A2 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__A2 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__A2 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__A2 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A2 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__A2 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__A2 (.I(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__I (.I(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__I (.I(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__I (.I(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A2 (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A2 (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A2 (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A2 (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__A2 (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A2 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A2 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A2 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__A2 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__A2 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A2 (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A2 (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__A2 (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A2 (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__A2 (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__A2 (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__I (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__I (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__I (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__A2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__A2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__A2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__A2 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A2 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__A2 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A2 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__A2 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__A2 (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__A2 (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__A2 (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__A2 (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__A2 (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11500__A2 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11489__I (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__I (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11483__I (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__A2 (.I(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__I (.I(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__I (.I(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__I (.I(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A2 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A2 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11534__A2 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__A2 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__A2 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__A2 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__I (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__I (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__I (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A2 (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__A2 (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A2 (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__A2 (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__A2 (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__A2 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__A2 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__A2 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A2 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11550__A2 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__C2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__A4 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__I (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__B (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__I (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__I (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__I1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A2 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__I0 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__I1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A2 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__I1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A2 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__I0 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__I1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A2 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__I1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__I1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A2 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__I1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A2 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A2 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A1 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A2 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__I0 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A2 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__A1 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__I0 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A1 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__A1 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A1 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A1 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A1 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A1 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A1 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__A1 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__I1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A2 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__I1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A2 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__I1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__I1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__A1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__I1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A2 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__I1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__I (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__I (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A2 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__B (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__I (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__S0 (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A1 (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A1 (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__I (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__A1 (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A1 (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A3 (.I(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__I (.I(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__A3 (.I(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__A1 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__I (.I(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__I (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__I (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__I (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__A2 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__I (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__I (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A3 (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A2 (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__A1 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__A1 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__B2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__I (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__B (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__I (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A2 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__B (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__I (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__B2 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A1 (.I(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__B2 (.I(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A2 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__C (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__I (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__B1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A2 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__I (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__B (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__C (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A2 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A2 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A2 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A2 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A1 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A2 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A1 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A1 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A1 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__I (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A1 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__B (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__A1 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__I (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05852__I (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__I (.I(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__I (.I(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__I (.I(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__A1 (.I(\u_cpu.rf_ram.memory[100][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__I0 (.I(\u_cpu.rf_ram.memory[100][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__A1 (.I(\u_cpu.rf_ram.memory[100][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__I0 (.I(\u_cpu.rf_ram.memory[100][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__A1 (.I(\u_cpu.rf_ram.memory[100][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__I0 (.I(\u_cpu.rf_ram.memory[100][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A1 (.I(\u_cpu.rf_ram.memory[100][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__I0 (.I(\u_cpu.rf_ram.memory[100][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__A1 (.I(\u_cpu.rf_ram.memory[100][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__I0 (.I(\u_cpu.rf_ram.memory[100][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A1 (.I(\u_cpu.rf_ram.memory[100][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__I0 (.I(\u_cpu.rf_ram.memory[100][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A1 (.I(\u_cpu.rf_ram.memory[100][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__I0 (.I(\u_cpu.rf_ram.memory[100][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(\u_cpu.rf_ram.memory[101][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__I1 (.I(\u_cpu.rf_ram.memory[101][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A1 (.I(\u_cpu.rf_ram.memory[101][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__I1 (.I(\u_cpu.rf_ram.memory[101][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A1 (.I(\u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__I2 (.I(\u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A1 (.I(\u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__I2 (.I(\u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(\u_cpu.rf_ram.memory[102][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__I2 (.I(\u_cpu.rf_ram.memory[102][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__A1 (.I(\u_cpu.rf_ram.memory[102][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__I2 (.I(\u_cpu.rf_ram.memory[102][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A1 (.I(\u_cpu.rf_ram.memory[102][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__I2 (.I(\u_cpu.rf_ram.memory[102][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(\u_cpu.rf_ram.memory[102][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__I2 (.I(\u_cpu.rf_ram.memory[102][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A1 (.I(\u_cpu.rf_ram.memory[103][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__I3 (.I(\u_cpu.rf_ram.memory[103][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A1 (.I(\u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__I0 (.I(\u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A1 (.I(\u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__I0 (.I(\u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A1 (.I(\u_cpu.rf_ram.memory[104][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__I0 (.I(\u_cpu.rf_ram.memory[104][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(\u_cpu.rf_ram.memory[106][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__I2 (.I(\u_cpu.rf_ram.memory[106][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A1 (.I(\u_cpu.rf_ram.memory[106][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__I2 (.I(\u_cpu.rf_ram.memory[106][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A1 (.I(\u_cpu.rf_ram.memory[106][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__I2 (.I(\u_cpu.rf_ram.memory[106][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A1 (.I(\u_cpu.rf_ram.memory[106][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__I2 (.I(\u_cpu.rf_ram.memory[106][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A1 (.I(\u_cpu.rf_ram.memory[106][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__I2 (.I(\u_cpu.rf_ram.memory[106][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(\u_cpu.rf_ram.memory[106][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__I2 (.I(\u_cpu.rf_ram.memory[106][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A1 (.I(\u_cpu.rf_ram.memory[106][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__I2 (.I(\u_cpu.rf_ram.memory[106][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A1 (.I(\u_cpu.rf_ram.memory[106][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__I2 (.I(\u_cpu.rf_ram.memory[106][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A1 (.I(\u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__I3 (.I(\u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A1 (.I(\u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__I3 (.I(\u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A1 (.I(\u_cpu.rf_ram.memory[107][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__I3 (.I(\u_cpu.rf_ram.memory[107][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__A1 (.I(\u_cpu.rf_ram.memory[107][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__I3 (.I(\u_cpu.rf_ram.memory[107][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__A1 (.I(\u_cpu.rf_ram.memory[107][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__I3 (.I(\u_cpu.rf_ram.memory[107][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__A1 (.I(\u_cpu.rf_ram.memory[107][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__I3 (.I(\u_cpu.rf_ram.memory[107][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__A1 (.I(\u_cpu.rf_ram.memory[107][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__I3 (.I(\u_cpu.rf_ram.memory[107][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A1 (.I(\u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I1 (.I(\u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A1 (.I(\u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__I1 (.I(\u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__A1 (.I(\u_cpu.rf_ram.memory[109][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I1 (.I(\u_cpu.rf_ram.memory[109][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__A1 (.I(\u_cpu.rf_ram.memory[109][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__I1 (.I(\u_cpu.rf_ram.memory[109][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(\u_cpu.rf_ram.memory[109][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__I1 (.I(\u_cpu.rf_ram.memory[109][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__A1 (.I(\u_cpu.rf_ram.memory[109][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__I1 (.I(\u_cpu.rf_ram.memory[109][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A1 (.I(\u_cpu.rf_ram.memory[109][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__I1 (.I(\u_cpu.rf_ram.memory[109][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__A1 (.I(\u_cpu.rf_ram.memory[109][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__I1 (.I(\u_cpu.rf_ram.memory[109][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A1 (.I(\u_cpu.rf_ram.memory[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__I2 (.I(\u_cpu.rf_ram.memory[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A1 (.I(\u_cpu.rf_ram.memory[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__I2 (.I(\u_cpu.rf_ram.memory[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A1 (.I(\u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I2 (.I(\u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__A1 (.I(\u_cpu.rf_ram.memory[110][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__I2 (.I(\u_cpu.rf_ram.memory[110][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A1 (.I(\u_cpu.rf_ram.memory[110][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I2 (.I(\u_cpu.rf_ram.memory[110][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A1 (.I(\u_cpu.rf_ram.memory[110][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__I2 (.I(\u_cpu.rf_ram.memory[110][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__A1 (.I(\u_cpu.rf_ram.memory[110][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__I2 (.I(\u_cpu.rf_ram.memory[110][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A1 (.I(\u_cpu.rf_ram.memory[110][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__I2 (.I(\u_cpu.rf_ram.memory[110][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A1 (.I(\u_cpu.rf_ram.memory[110][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__I2 (.I(\u_cpu.rf_ram.memory[110][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A1 (.I(\u_cpu.rf_ram.memory[110][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__I2 (.I(\u_cpu.rf_ram.memory[110][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(\u_cpu.rf_ram.memory[111][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I3 (.I(\u_cpu.rf_ram.memory[111][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__A1 (.I(\u_cpu.rf_ram.memory[111][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__I3 (.I(\u_cpu.rf_ram.memory[111][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(\u_cpu.rf_ram.memory[111][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I3 (.I(\u_cpu.rf_ram.memory[111][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A1 (.I(\u_cpu.rf_ram.memory[112][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__I0 (.I(\u_cpu.rf_ram.memory[112][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A1 (.I(\u_cpu.rf_ram.memory[112][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__I0 (.I(\u_cpu.rf_ram.memory[112][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(\u_cpu.rf_ram.memory[112][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__I0 (.I(\u_cpu.rf_ram.memory[112][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A1 (.I(\u_cpu.rf_ram.memory[112][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__I0 (.I(\u_cpu.rf_ram.memory[112][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A1 (.I(\u_cpu.rf_ram.memory[112][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__I0 (.I(\u_cpu.rf_ram.memory[112][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__A1 (.I(\u_cpu.rf_ram.memory[114][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__I2 (.I(\u_cpu.rf_ram.memory[114][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A1 (.I(\u_cpu.rf_ram.memory[114][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__I2 (.I(\u_cpu.rf_ram.memory[114][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A1 (.I(\u_cpu.rf_ram.memory[114][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__I2 (.I(\u_cpu.rf_ram.memory[114][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(\u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__I0 (.I(\u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(\u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I0 (.I(\u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(\u_cpu.rf_ram.memory[116][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__I0 (.I(\u_cpu.rf_ram.memory[116][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(\u_cpu.rf_ram.memory[116][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__I0 (.I(\u_cpu.rf_ram.memory[116][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A1 (.I(\u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I1 (.I(\u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A1 (.I(\u_cpu.rf_ram.memory[117][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__I1 (.I(\u_cpu.rf_ram.memory[117][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A1 (.I(\u_cpu.rf_ram.memory[117][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__I1 (.I(\u_cpu.rf_ram.memory[117][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(\u_cpu.rf_ram.memory[117][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__I1 (.I(\u_cpu.rf_ram.memory[117][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(\u_cpu.rf_ram.memory[117][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__I1 (.I(\u_cpu.rf_ram.memory[117][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(\u_cpu.rf_ram.memory[118][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__I2 (.I(\u_cpu.rf_ram.memory[118][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A1 (.I(\u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__I3 (.I(\u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A1 (.I(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I3 (.I(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A1 (.I(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__I3 (.I(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A1 (.I(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__I3 (.I(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__I3 (.I(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A1 (.I(\u_cpu.rf_ram.memory[119][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__I3 (.I(\u_cpu.rf_ram.memory[119][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A1 (.I(\u_cpu.rf_ram.memory[119][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__I3 (.I(\u_cpu.rf_ram.memory[119][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A1 (.I(\u_cpu.rf_ram.memory[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__I3 (.I(\u_cpu.rf_ram.memory[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A1 (.I(\u_cpu.rf_ram.memory[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__I3 (.I(\u_cpu.rf_ram.memory[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(\u_cpu.rf_ram.memory[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__I3 (.I(\u_cpu.rf_ram.memory[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(\u_cpu.rf_ram.memory[120][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__I0 (.I(\u_cpu.rf_ram.memory[120][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(\u_cpu.rf_ram.memory[120][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__I0 (.I(\u_cpu.rf_ram.memory[120][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(\u_cpu.rf_ram.memory[120][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__I0 (.I(\u_cpu.rf_ram.memory[120][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(\u_cpu.rf_ram.memory[120][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__I0 (.I(\u_cpu.rf_ram.memory[120][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__I0 (.I(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A1 (.I(\u_cpu.rf_ram.memory[120][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__I0 (.I(\u_cpu.rf_ram.memory[120][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A1 (.I(\u_cpu.rf_ram.memory[120][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__I0 (.I(\u_cpu.rf_ram.memory[120][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A1 (.I(\u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__I2 (.I(\u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(\u_cpu.rf_ram.memory[122][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__I2 (.I(\u_cpu.rf_ram.memory[122][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A1 (.I(\u_cpu.rf_ram.memory[122][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__I2 (.I(\u_cpu.rf_ram.memory[122][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A1 (.I(\u_cpu.rf_ram.memory[123][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__I3 (.I(\u_cpu.rf_ram.memory[123][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A1 (.I(\u_cpu.rf_ram.memory[123][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__I3 (.I(\u_cpu.rf_ram.memory[123][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A1 (.I(\u_cpu.rf_ram.memory[124][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__I0 (.I(\u_cpu.rf_ram.memory[124][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A1 (.I(\u_cpu.rf_ram.memory[124][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__I0 (.I(\u_cpu.rf_ram.memory[124][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A1 (.I(\u_cpu.rf_ram.memory[124][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__I0 (.I(\u_cpu.rf_ram.memory[124][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A1 (.I(\u_cpu.rf_ram.memory[124][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__I0 (.I(\u_cpu.rf_ram.memory[124][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A1 (.I(\u_cpu.rf_ram.memory[124][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__I0 (.I(\u_cpu.rf_ram.memory[124][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A1 (.I(\u_cpu.rf_ram.memory[124][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__I0 (.I(\u_cpu.rf_ram.memory[124][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__I0 (.I(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A1 (.I(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__I0 (.I(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A1 (.I(\u_cpu.rf_ram.memory[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__I0 (.I(\u_cpu.rf_ram.memory[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A1 (.I(\u_cpu.rf_ram.memory[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I0 (.I(\u_cpu.rf_ram.memory[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A1 (.I(\u_cpu.rf_ram.memory[128][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__I0 (.I(\u_cpu.rf_ram.memory[128][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A1 (.I(\u_cpu.rf_ram.memory[128][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__I0 (.I(\u_cpu.rf_ram.memory[128][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A1 (.I(\u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__I1 (.I(\u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(\u_cpu.rf_ram.memory[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__I1 (.I(\u_cpu.rf_ram.memory[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A1 (.I(\u_cpu.rf_ram.memory[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__I1 (.I(\u_cpu.rf_ram.memory[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A1 (.I(\u_cpu.rf_ram.memory[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__I1 (.I(\u_cpu.rf_ram.memory[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(\u_cpu.rf_ram.memory[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__I0 (.I(\u_cpu.rf_ram.memory[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(\u_cpu.rf_ram.memory[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__I0 (.I(\u_cpu.rf_ram.memory[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A1 (.I(\u_cpu.rf_ram.memory[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__I0 (.I(\u_cpu.rf_ram.memory[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(\u_cpu.rf_ram.memory[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__I0 (.I(\u_cpu.rf_ram.memory[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A1 (.I(\u_cpu.rf_ram.memory[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__I0 (.I(\u_cpu.rf_ram.memory[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A1 (.I(\u_cpu.rf_ram.memory[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__I0 (.I(\u_cpu.rf_ram.memory[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(\u_cpu.rf_ram.memory[130][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__I2 (.I(\u_cpu.rf_ram.memory[130][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(\u_cpu.rf_ram.memory[131][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__I3 (.I(\u_cpu.rf_ram.memory[131][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(\u_cpu.rf_ram.memory[131][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__I3 (.I(\u_cpu.rf_ram.memory[131][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(\u_cpu.rf_ram.memory[135][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__I3 (.I(\u_cpu.rf_ram.memory[135][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(\u_cpu.rf_ram.memory[135][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__I3 (.I(\u_cpu.rf_ram.memory[135][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(\u_cpu.rf_ram.memory[135][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__I3 (.I(\u_cpu.rf_ram.memory[135][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A1 (.I(\u_cpu.rf_ram.memory[135][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__I3 (.I(\u_cpu.rf_ram.memory[135][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(\u_cpu.rf_ram.memory[135][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__I3 (.I(\u_cpu.rf_ram.memory[135][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A1 (.I(\u_cpu.rf_ram.memory[135][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__I3 (.I(\u_cpu.rf_ram.memory[135][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A1 (.I(\u_cpu.rf_ram.memory[135][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__I3 (.I(\u_cpu.rf_ram.memory[135][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A1 (.I(\u_cpu.rf_ram.memory[135][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__I3 (.I(\u_cpu.rf_ram.memory[135][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A1 (.I(\u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__I0 (.I(\u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A1 (.I(\u_cpu.rf_ram.memory[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__I0 (.I(\u_cpu.rf_ram.memory[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A1 (.I(\u_cpu.rf_ram.memory[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__I0 (.I(\u_cpu.rf_ram.memory[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A1 (.I(\u_cpu.rf_ram.memory[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I0 (.I(\u_cpu.rf_ram.memory[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A1 (.I(\u_cpu.rf_ram.memory[136][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__I0 (.I(\u_cpu.rf_ram.memory[136][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A1 (.I(\u_cpu.rf_ram.memory[136][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__I0 (.I(\u_cpu.rf_ram.memory[136][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A1 (.I(\u_cpu.rf_ram.memory[137][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__I1 (.I(\u_cpu.rf_ram.memory[137][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A1 (.I(\u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__I2 (.I(\u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A1 (.I(\u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__I2 (.I(\u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A1 (.I(\u_cpu.rf_ram.memory[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__I2 (.I(\u_cpu.rf_ram.memory[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A1 (.I(\u_cpu.rf_ram.memory[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__I2 (.I(\u_cpu.rf_ram.memory[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(\u_cpu.rf_ram.memory[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I2 (.I(\u_cpu.rf_ram.memory[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__A1 (.I(\u_cpu.rf_ram.memory[138][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__I2 (.I(\u_cpu.rf_ram.memory[138][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A1 (.I(\u_cpu.rf_ram.memory[138][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__I2 (.I(\u_cpu.rf_ram.memory[138][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(\u_cpu.rf_ram.memory[138][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__I2 (.I(\u_cpu.rf_ram.memory[138][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A1 (.I(\u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__I3 (.I(\u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A1 (.I(\u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__I3 (.I(\u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A1 (.I(\u_cpu.rf_ram.memory[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__I3 (.I(\u_cpu.rf_ram.memory[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A1 (.I(\u_cpu.rf_ram.memory[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__I3 (.I(\u_cpu.rf_ram.memory[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A1 (.I(\u_cpu.rf_ram.memory[139][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I3 (.I(\u_cpu.rf_ram.memory[139][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A1 (.I(\u_cpu.rf_ram.memory[139][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__I3 (.I(\u_cpu.rf_ram.memory[139][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A1 (.I(\u_cpu.rf_ram.memory[142][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__I2 (.I(\u_cpu.rf_ram.memory[142][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(\u_cpu.rf_ram.memory[142][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__I2 (.I(\u_cpu.rf_ram.memory[142][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(\u_cpu.rf_ram.memory[142][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__I2 (.I(\u_cpu.rf_ram.memory[142][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(\u_cpu.rf_ram.memory[143][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__I3 (.I(\u_cpu.rf_ram.memory[143][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(\u_cpu.rf_ram.memory[143][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__I3 (.I(\u_cpu.rf_ram.memory[143][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(\u_cpu.rf_ram.memory[143][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__I3 (.I(\u_cpu.rf_ram.memory[143][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(\u_cpu.rf_ram.memory[143][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__I3 (.I(\u_cpu.rf_ram.memory[143][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A1 (.I(\u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__I2 (.I(\u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(\u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__I2 (.I(\u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A1 (.I(\u_cpu.rf_ram.memory[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__I2 (.I(\u_cpu.rf_ram.memory[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(\u_cpu.rf_ram.memory[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__I2 (.I(\u_cpu.rf_ram.memory[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(\u_cpu.rf_ram.memory[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__I2 (.I(\u_cpu.rf_ram.memory[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(\u_cpu.rf_ram.memory[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__I2 (.I(\u_cpu.rf_ram.memory[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A1 (.I(\u_cpu.rf_ram.memory[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__I2 (.I(\u_cpu.rf_ram.memory[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(\u_cpu.rf_ram.memory[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__I2 (.I(\u_cpu.rf_ram.memory[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A1 (.I(\u_cpu.rf_ram.memory[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__I3 (.I(\u_cpu.rf_ram.memory[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A1 (.I(\u_cpu.rf_ram.memory[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__I0 (.I(\u_cpu.rf_ram.memory[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A1 (.I(\u_cpu.rf_ram.memory[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__I0 (.I(\u_cpu.rf_ram.memory[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A1 (.I(\u_cpu.rf_ram.memory[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__I0 (.I(\u_cpu.rf_ram.memory[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A1 (.I(\u_cpu.rf_ram.memory[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__I0 (.I(\u_cpu.rf_ram.memory[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A1 (.I(\u_cpu.rf_ram.memory[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__I0 (.I(\u_cpu.rf_ram.memory[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A1 (.I(\u_cpu.rf_ram.memory[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__I0 (.I(\u_cpu.rf_ram.memory[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A1 (.I(\u_cpu.rf_ram.memory[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__I0 (.I(\u_cpu.rf_ram.memory[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A1 (.I(\u_cpu.rf_ram.memory[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__I0 (.I(\u_cpu.rf_ram.memory[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A1 (.I(\u_cpu.rf_ram.memory[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__I1 (.I(\u_cpu.rf_ram.memory[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A1 (.I(\u_cpu.rf_ram.memory[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__I1 (.I(\u_cpu.rf_ram.memory[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A1 (.I(\u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__I3 (.I(\u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A1 (.I(\u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__I3 (.I(\u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__I3 (.I(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A1 (.I(\u_cpu.rf_ram.memory[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__I3 (.I(\u_cpu.rf_ram.memory[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A1 (.I(\u_cpu.rf_ram.memory[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__I3 (.I(\u_cpu.rf_ram.memory[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A1 (.I(\u_cpu.rf_ram.memory[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__I3 (.I(\u_cpu.rf_ram.memory[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A1 (.I(\u_cpu.rf_ram.memory[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__I3 (.I(\u_cpu.rf_ram.memory[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__I3 (.I(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A1 (.I(\u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__I1 (.I(\u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(\u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__I1 (.I(\u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A1 (.I(\u_cpu.rf_ram.memory[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__I1 (.I(\u_cpu.rf_ram.memory[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(\u_cpu.rf_ram.memory[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__I1 (.I(\u_cpu.rf_ram.memory[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A1 (.I(\u_cpu.rf_ram.memory[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__I1 (.I(\u_cpu.rf_ram.memory[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A1 (.I(\u_cpu.rf_ram.memory[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__I1 (.I(\u_cpu.rf_ram.memory[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A1 (.I(\u_cpu.rf_ram.memory[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__I1 (.I(\u_cpu.rf_ram.memory[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A1 (.I(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__I2 (.I(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__I2 (.I(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(\u_cpu.rf_ram.memory[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__I2 (.I(\u_cpu.rf_ram.memory[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A1 (.I(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__I2 (.I(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A1 (.I(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__I2 (.I(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A1 (.I(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__I2 (.I(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A1 (.I(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__I2 (.I(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__I2 (.I(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11550__A1 (.I(\u_cpu.rf_ram.memory[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__I3 (.I(\u_cpu.rf_ram.memory[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A1 (.I(\u_cpu.rf_ram.memory[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__I3 (.I(\u_cpu.rf_ram.memory[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__A1 (.I(\u_cpu.rf_ram.memory[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__I3 (.I(\u_cpu.rf_ram.memory[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__A1 (.I(\u_cpu.rf_ram.memory[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__I3 (.I(\u_cpu.rf_ram.memory[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A1 (.I(\u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__I0 (.I(\u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A1 (.I(\u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__I0 (.I(\u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A1 (.I(\u_cpu.rf_ram.memory[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__I0 (.I(\u_cpu.rf_ram.memory[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__A1 (.I(\u_cpu.rf_ram.memory[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__I0 (.I(\u_cpu.rf_ram.memory[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A1 (.I(\u_cpu.rf_ram.memory[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__I0 (.I(\u_cpu.rf_ram.memory[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A1 (.I(\u_cpu.rf_ram.memory[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__I0 (.I(\u_cpu.rf_ram.memory[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A1 (.I(\u_cpu.rf_ram.memory[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__I0 (.I(\u_cpu.rf_ram.memory[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__A1 (.I(\u_cpu.rf_ram.memory[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__I0 (.I(\u_cpu.rf_ram.memory[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__I1 (.I(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A1 (.I(\u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__I1 (.I(\u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__A1 (.I(\u_cpu.rf_ram.memory[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__I1 (.I(\u_cpu.rf_ram.memory[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(\u_cpu.rf_ram.memory[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__I1 (.I(\u_cpu.rf_ram.memory[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A1 (.I(\u_cpu.rf_ram.memory[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__I2 (.I(\u_cpu.rf_ram.memory[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A1 (.I(\u_cpu.rf_ram.memory[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__I2 (.I(\u_cpu.rf_ram.memory[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A1 (.I(\u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__I0 (.I(\u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A1 (.I(\u_cpu.rf_ram.memory[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__I0 (.I(\u_cpu.rf_ram.memory[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A1 (.I(\u_cpu.rf_ram.memory[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I0 (.I(\u_cpu.rf_ram.memory[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__A1 (.I(\u_cpu.rf_ram.memory[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__I0 (.I(\u_cpu.rf_ram.memory[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(\u_cpu.rf_ram.memory[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__I0 (.I(\u_cpu.rf_ram.memory[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(\u_cpu.rf_ram.memory[33][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__I1 (.I(\u_cpu.rf_ram.memory[33][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A1 (.I(\u_cpu.rf_ram.memory[33][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__I1 (.I(\u_cpu.rf_ram.memory[33][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(\u_cpu.rf_ram.memory[35][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__I3 (.I(\u_cpu.rf_ram.memory[35][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A1 (.I(\u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__I0 (.I(\u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A1 (.I(\u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__I0 (.I(\u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__A1 (.I(\u_cpu.rf_ram.memory[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__I0 (.I(\u_cpu.rf_ram.memory[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A1 (.I(\u_cpu.rf_ram.memory[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__I0 (.I(\u_cpu.rf_ram.memory[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(\u_cpu.rf_ram.memory[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__I0 (.I(\u_cpu.rf_ram.memory[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A1 (.I(\u_cpu.rf_ram.memory[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__I0 (.I(\u_cpu.rf_ram.memory[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A1 (.I(\u_cpu.rf_ram.memory[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__I0 (.I(\u_cpu.rf_ram.memory[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(\u_cpu.rf_ram.memory[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__I1 (.I(\u_cpu.rf_ram.memory[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A1 (.I(\u_cpu.rf_ram.memory[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__I1 (.I(\u_cpu.rf_ram.memory[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A1 (.I(\u_cpu.rf_ram.memory[37][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__I1 (.I(\u_cpu.rf_ram.memory[37][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A1 (.I(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__I3 (.I(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__I3 (.I(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__I3 (.I(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(\u_cpu.rf_ram.memory[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__I3 (.I(\u_cpu.rf_ram.memory[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A1 (.I(\u_cpu.rf_ram.memory[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__I3 (.I(\u_cpu.rf_ram.memory[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__I3 (.I(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(\u_cpu.rf_ram.memory[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__I3 (.I(\u_cpu.rf_ram.memory[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A1 (.I(\u_cpu.rf_ram.memory[40][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__I0 (.I(\u_cpu.rf_ram.memory[40][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A1 (.I(\u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__I1 (.I(\u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A1 (.I(\u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__I1 (.I(\u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A1 (.I(\u_cpu.rf_ram.memory[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__I1 (.I(\u_cpu.rf_ram.memory[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(\u_cpu.rf_ram.memory[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__I1 (.I(\u_cpu.rf_ram.memory[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A1 (.I(\u_cpu.rf_ram.memory[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__I1 (.I(\u_cpu.rf_ram.memory[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A1 (.I(\u_cpu.rf_ram.memory[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__I1 (.I(\u_cpu.rf_ram.memory[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A1 (.I(\u_cpu.rf_ram.memory[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__I1 (.I(\u_cpu.rf_ram.memory[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A1 (.I(\u_cpu.rf_ram.memory[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__I1 (.I(\u_cpu.rf_ram.memory[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A1 (.I(\u_cpu.rf_ram.memory[42][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__I2 (.I(\u_cpu.rf_ram.memory[42][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A1 (.I(\u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__I0 (.I(\u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A1 (.I(\u_cpu.rf_ram.memory[44][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__I0 (.I(\u_cpu.rf_ram.memory[44][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A1 (.I(\u_cpu.rf_ram.memory[44][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__I0 (.I(\u_cpu.rf_ram.memory[44][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__A1 (.I(\u_cpu.rf_ram.memory[44][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__I0 (.I(\u_cpu.rf_ram.memory[44][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A1 (.I(\u_cpu.rf_ram.memory[44][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__I0 (.I(\u_cpu.rf_ram.memory[44][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A1 (.I(\u_cpu.rf_ram.memory[44][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__I0 (.I(\u_cpu.rf_ram.memory[44][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A1 (.I(\u_cpu.rf_ram.memory[45][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__I1 (.I(\u_cpu.rf_ram.memory[45][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A1 (.I(\u_cpu.rf_ram.memory[45][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__I1 (.I(\u_cpu.rf_ram.memory[45][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__A1 (.I(\u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__I2 (.I(\u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__A1 (.I(\u_cpu.rf_ram.memory[46][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__I2 (.I(\u_cpu.rf_ram.memory[46][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__A1 (.I(\u_cpu.rf_ram.memory[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__I2 (.I(\u_cpu.rf_ram.memory[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A1 (.I(\u_cpu.rf_ram.memory[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__I2 (.I(\u_cpu.rf_ram.memory[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A1 (.I(\u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__I3 (.I(\u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__A1 (.I(\u_cpu.rf_ram.memory[48][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__I0 (.I(\u_cpu.rf_ram.memory[48][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__I1 (.I(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__I1 (.I(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A1 (.I(\u_cpu.rf_ram.memory[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__I1 (.I(\u_cpu.rf_ram.memory[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A1 (.I(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__I1 (.I(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A1 (.I(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__I1 (.I(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__I1 (.I(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A1 (.I(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__I1 (.I(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(\u_cpu.rf_ram.memory[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__I1 (.I(\u_cpu.rf_ram.memory[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A1 (.I(\u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__I3 (.I(\u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__A1 (.I(\u_cpu.rf_ram.memory[51][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__I3 (.I(\u_cpu.rf_ram.memory[51][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A1 (.I(\u_cpu.rf_ram.memory[51][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__I3 (.I(\u_cpu.rf_ram.memory[51][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A1 (.I(\u_cpu.rf_ram.memory[51][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__I3 (.I(\u_cpu.rf_ram.memory[51][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__A1 (.I(\u_cpu.rf_ram.memory[51][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__I3 (.I(\u_cpu.rf_ram.memory[51][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(\u_cpu.rf_ram.memory[52][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__I0 (.I(\u_cpu.rf_ram.memory[52][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A1 (.I(\u_cpu.rf_ram.memory[54][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__I2 (.I(\u_cpu.rf_ram.memory[54][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A1 (.I(\u_cpu.rf_ram.memory[54][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__I2 (.I(\u_cpu.rf_ram.memory[54][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(\u_cpu.rf_ram.memory[54][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__I2 (.I(\u_cpu.rf_ram.memory[54][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(\u_cpu.rf_ram.memory[54][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__I2 (.I(\u_cpu.rf_ram.memory[54][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(\u_cpu.rf_ram.memory[54][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__I2 (.I(\u_cpu.rf_ram.memory[54][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A1 (.I(\u_cpu.rf_ram.memory[54][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__I2 (.I(\u_cpu.rf_ram.memory[54][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(\u_cpu.rf_ram.memory[55][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__I3 (.I(\u_cpu.rf_ram.memory[55][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A1 (.I(\u_cpu.rf_ram.memory[55][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__I3 (.I(\u_cpu.rf_ram.memory[55][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A1 (.I(\u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__I0 (.I(\u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A1 (.I(\u_cpu.rf_ram.memory[58][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__I2 (.I(\u_cpu.rf_ram.memory[58][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A1 (.I(\u_cpu.rf_ram.memory[58][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__I2 (.I(\u_cpu.rf_ram.memory[58][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A1 (.I(\u_cpu.rf_ram.memory[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__I2 (.I(\u_cpu.rf_ram.memory[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A1 (.I(\u_cpu.rf_ram.memory[58][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__I2 (.I(\u_cpu.rf_ram.memory[58][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(\u_cpu.rf_ram.memory[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__I2 (.I(\u_cpu.rf_ram.memory[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A1 (.I(\u_cpu.rf_ram.memory[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__I2 (.I(\u_cpu.rf_ram.memory[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(\u_cpu.rf_ram.memory[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__I2 (.I(\u_cpu.rf_ram.memory[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A1 (.I(\u_cpu.rf_ram.memory[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__I2 (.I(\u_cpu.rf_ram.memory[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A1 (.I(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__I3 (.I(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(\u_cpu.rf_ram.memory[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__I1 (.I(\u_cpu.rf_ram.memory[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A1 (.I(\u_cpu.rf_ram.memory[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__I1 (.I(\u_cpu.rf_ram.memory[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A1 (.I(\u_cpu.rf_ram.memory[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__I1 (.I(\u_cpu.rf_ram.memory[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A1 (.I(\u_cpu.rf_ram.memory[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__I1 (.I(\u_cpu.rf_ram.memory[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A1 (.I(\u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__I0 (.I(\u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A1 (.I(\u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__I0 (.I(\u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A1 (.I(\u_cpu.rf_ram.memory[60][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__I0 (.I(\u_cpu.rf_ram.memory[60][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A1 (.I(\u_cpu.rf_ram.memory[63][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__I3 (.I(\u_cpu.rf_ram.memory[63][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A1 (.I(\u_cpu.rf_ram.memory[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__I3 (.I(\u_cpu.rf_ram.memory[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A1 (.I(\u_cpu.rf_ram.memory[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__I3 (.I(\u_cpu.rf_ram.memory[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A1 (.I(\u_cpu.rf_ram.memory[63][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__I3 (.I(\u_cpu.rf_ram.memory[63][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A1 (.I(\u_cpu.rf_ram.memory[63][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__I3 (.I(\u_cpu.rf_ram.memory[63][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A1 (.I(\u_cpu.rf_ram.memory[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__I3 (.I(\u_cpu.rf_ram.memory[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A1 (.I(\u_cpu.rf_ram.memory[67][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__I3 (.I(\u_cpu.rf_ram.memory[67][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A1 (.I(\u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__I2 (.I(\u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(\u_cpu.rf_ram.memory[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__I2 (.I(\u_cpu.rf_ram.memory[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(\u_cpu.rf_ram.memory[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__I2 (.I(\u_cpu.rf_ram.memory[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A1 (.I(\u_cpu.rf_ram.memory[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__I2 (.I(\u_cpu.rf_ram.memory[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A1 (.I(\u_cpu.rf_ram.memory[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__I2 (.I(\u_cpu.rf_ram.memory[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A1 (.I(\u_cpu.rf_ram.memory[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__I2 (.I(\u_cpu.rf_ram.memory[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A1 (.I(\u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__I2 (.I(\u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A1 (.I(\u_cpu.rf_ram.memory[70][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__I2 (.I(\u_cpu.rf_ram.memory[70][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A1 (.I(\u_cpu.rf_ram.memory[70][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__I2 (.I(\u_cpu.rf_ram.memory[70][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A1 (.I(\u_cpu.rf_ram.memory[70][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__I2 (.I(\u_cpu.rf_ram.memory[70][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(\u_cpu.rf_ram.memory[70][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__I2 (.I(\u_cpu.rf_ram.memory[70][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A1 (.I(\u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__I3 (.I(\u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(\u_cpu.rf_ram.memory[71][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__I3 (.I(\u_cpu.rf_ram.memory[71][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(\u_cpu.rf_ram.memory[71][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__I3 (.I(\u_cpu.rf_ram.memory[71][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__A1 (.I(\u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__I0 (.I(\u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(\u_cpu.rf_ram.memory[72][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__I0 (.I(\u_cpu.rf_ram.memory[72][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A1 (.I(\u_cpu.rf_ram.memory[72][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__I0 (.I(\u_cpu.rf_ram.memory[72][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A1 (.I(\u_cpu.rf_ram.memory[72][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__I0 (.I(\u_cpu.rf_ram.memory[72][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A1 (.I(\u_cpu.rf_ram.memory[72][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__I0 (.I(\u_cpu.rf_ram.memory[72][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(\u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__I1 (.I(\u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(\u_cpu.rf_ram.memory[73][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__I1 (.I(\u_cpu.rf_ram.memory[73][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(\u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__I0 (.I(\u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A1 (.I(\u_cpu.rf_ram.memory[76][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__I0 (.I(\u_cpu.rf_ram.memory[76][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(\u_cpu.rf_ram.memory[77][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__I1 (.I(\u_cpu.rf_ram.memory[77][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A1 (.I(\u_cpu.rf_ram.memory[77][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__I1 (.I(\u_cpu.rf_ram.memory[77][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(\u_cpu.rf_ram.memory[77][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__I1 (.I(\u_cpu.rf_ram.memory[77][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(\u_cpu.rf_ram.memory[77][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I1 (.I(\u_cpu.rf_ram.memory[77][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A1 (.I(\u_cpu.rf_ram.memory[77][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__I1 (.I(\u_cpu.rf_ram.memory[77][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A1 (.I(\u_cpu.rf_ram.memory[77][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__I1 (.I(\u_cpu.rf_ram.memory[77][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(\u_cpu.rf_ram.memory[77][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__I1 (.I(\u_cpu.rf_ram.memory[77][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A1 (.I(\u_cpu.rf_ram.memory[77][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__I1 (.I(\u_cpu.rf_ram.memory[77][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A1 (.I(\u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__I2 (.I(\u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__A1 (.I(\u_cpu.rf_ram.memory[78][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__I2 (.I(\u_cpu.rf_ram.memory[78][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__A1 (.I(\u_cpu.rf_ram.memory[78][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I2 (.I(\u_cpu.rf_ram.memory[78][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A1 (.I(\u_cpu.rf_ram.memory[78][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__I2 (.I(\u_cpu.rf_ram.memory[78][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A1 (.I(\u_cpu.rf_ram.memory[78][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__I2 (.I(\u_cpu.rf_ram.memory[78][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A1 (.I(\u_cpu.rf_ram.memory[78][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__I2 (.I(\u_cpu.rf_ram.memory[78][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A1 (.I(\u_cpu.rf_ram.memory[78][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__I2 (.I(\u_cpu.rf_ram.memory[78][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A1 (.I(\u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__I3 (.I(\u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A1 (.I(\u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__I3 (.I(\u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__A1 (.I(\u_cpu.rf_ram.memory[79][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__I3 (.I(\u_cpu.rf_ram.memory[79][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__A1 (.I(\u_cpu.rf_ram.memory[79][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I3 (.I(\u_cpu.rf_ram.memory[79][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A1 (.I(\u_cpu.rf_ram.memory[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__I3 (.I(\u_cpu.rf_ram.memory[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A1 (.I(\u_cpu.rf_ram.memory[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__I3 (.I(\u_cpu.rf_ram.memory[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A1 (.I(\u_cpu.rf_ram.memory[81][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I1 (.I(\u_cpu.rf_ram.memory[81][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(\u_cpu.rf_ram.memory[81][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__I1 (.I(\u_cpu.rf_ram.memory[81][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A1 (.I(\u_cpu.rf_ram.memory[81][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__I1 (.I(\u_cpu.rf_ram.memory[81][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A1 (.I(\u_cpu.rf_ram.memory[81][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__I1 (.I(\u_cpu.rf_ram.memory[81][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A1 (.I(\u_cpu.rf_ram.memory[81][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__I1 (.I(\u_cpu.rf_ram.memory[81][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A1 (.I(\u_cpu.rf_ram.memory[81][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__I1 (.I(\u_cpu.rf_ram.memory[81][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__A1 (.I(\u_cpu.rf_ram.memory[82][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I2 (.I(\u_cpu.rf_ram.memory[82][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A1 (.I(\u_cpu.rf_ram.memory[82][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__I2 (.I(\u_cpu.rf_ram.memory[82][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(\u_cpu.rf_ram.memory[82][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__I2 (.I(\u_cpu.rf_ram.memory[82][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(\u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__I3 (.I(\u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A1 (.I(\u_cpu.rf_ram.memory[83][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__I3 (.I(\u_cpu.rf_ram.memory[83][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A1 (.I(\u_cpu.rf_ram.memory[83][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__I3 (.I(\u_cpu.rf_ram.memory[83][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A1 (.I(\u_cpu.rf_ram.memory[83][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__I3 (.I(\u_cpu.rf_ram.memory[83][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A1 (.I(\u_cpu.rf_ram.memory[83][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__I3 (.I(\u_cpu.rf_ram.memory[83][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__A1 (.I(\u_cpu.rf_ram.memory[84][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__I0 (.I(\u_cpu.rf_ram.memory[84][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__A1 (.I(\u_cpu.rf_ram.memory[84][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__I0 (.I(\u_cpu.rf_ram.memory[84][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A1 (.I(\u_cpu.rf_ram.memory[88][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__I0 (.I(\u_cpu.rf_ram.memory[88][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(\u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__I0 (.I(\u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A1 (.I(\u_cpu.rf_ram.memory[88][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__I0 (.I(\u_cpu.rf_ram.memory[88][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A1 (.I(\u_cpu.rf_ram.memory[88][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__I0 (.I(\u_cpu.rf_ram.memory[88][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__A1 (.I(\u_cpu.rf_ram.memory[88][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__I0 (.I(\u_cpu.rf_ram.memory[88][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(\u_cpu.rf_ram.memory[88][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__I0 (.I(\u_cpu.rf_ram.memory[88][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__A1 (.I(\u_cpu.rf_ram.memory[88][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__I0 (.I(\u_cpu.rf_ram.memory[88][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(\u_cpu.rf_ram.memory[88][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__I0 (.I(\u_cpu.rf_ram.memory[88][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__A1 (.I(\u_cpu.rf_ram.memory[89][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__I1 (.I(\u_cpu.rf_ram.memory[89][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11527__A1 (.I(\u_cpu.rf_ram.memory[89][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__I1 (.I(\u_cpu.rf_ram.memory[89][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__A1 (.I(\u_cpu.rf_ram.memory[89][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__I1 (.I(\u_cpu.rf_ram.memory[89][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__A1 (.I(\u_cpu.rf_ram.memory[89][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__I1 (.I(\u_cpu.rf_ram.memory[89][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11534__A1 (.I(\u_cpu.rf_ram.memory[89][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__I1 (.I(\u_cpu.rf_ram.memory[89][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A1 (.I(\u_cpu.rf_ram.memory[89][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__I1 (.I(\u_cpu.rf_ram.memory[89][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A1 (.I(\u_cpu.rf_ram.memory[89][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__I1 (.I(\u_cpu.rf_ram.memory[89][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11540__A1 (.I(\u_cpu.rf_ram.memory[89][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__I1 (.I(\u_cpu.rf_ram.memory[89][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(\u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__I0 (.I(\u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A1 (.I(\u_cpu.rf_ram.memory[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__I0 (.I(\u_cpu.rf_ram.memory[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(\u_cpu.rf_ram.memory[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__I0 (.I(\u_cpu.rf_ram.memory[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(\u_cpu.rf_ram.memory[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__I0 (.I(\u_cpu.rf_ram.memory[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A1 (.I(\u_cpu.rf_ram.memory[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__I0 (.I(\u_cpu.rf_ram.memory[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A1 (.I(\u_cpu.rf_ram.memory[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__I0 (.I(\u_cpu.rf_ram.memory[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(\u_cpu.rf_ram.memory[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__I0 (.I(\u_cpu.rf_ram.memory[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A1 (.I(\u_cpu.rf_ram.memory[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__I0 (.I(\u_cpu.rf_ram.memory[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A1 (.I(\u_cpu.rf_ram.memory[91][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__I3 (.I(\u_cpu.rf_ram.memory[91][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(\u_cpu.rf_ram.memory[91][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__I3 (.I(\u_cpu.rf_ram.memory[91][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A1 (.I(\u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__I0 (.I(\u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A1 (.I(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I0 (.I(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__I0 (.I(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(\u_cpu.rf_ram.memory[92][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__I0 (.I(\u_cpu.rf_ram.memory[92][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(\u_cpu.rf_ram.memory[92][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__I0 (.I(\u_cpu.rf_ram.memory[92][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A1 (.I(\u_cpu.rf_ram.memory[92][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__I0 (.I(\u_cpu.rf_ram.memory[92][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(\u_cpu.rf_ram.memory[92][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__I0 (.I(\u_cpu.rf_ram.memory[92][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A1 (.I(\u_cpu.rf_ram.memory[92][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__I0 (.I(\u_cpu.rf_ram.memory[92][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A1 (.I(\u_cpu.rf_ram.memory[94][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__I2 (.I(\u_cpu.rf_ram.memory[94][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A1 (.I(\u_cpu.rf_ram.memory[94][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__I2 (.I(\u_cpu.rf_ram.memory[94][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A1 (.I(\u_cpu.rf_ram.memory[94][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__I2 (.I(\u_cpu.rf_ram.memory[94][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A1 (.I(\u_cpu.rf_ram.memory[95][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I3 (.I(\u_cpu.rf_ram.memory[95][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A1 (.I(\u_cpu.rf_ram.memory[95][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__I3 (.I(\u_cpu.rf_ram.memory[95][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__A1 (.I(\u_cpu.rf_ram.memory[95][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__I3 (.I(\u_cpu.rf_ram.memory[95][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A1 (.I(\u_cpu.rf_ram.memory[95][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__I3 (.I(\u_cpu.rf_ram.memory[95][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A1 (.I(\u_cpu.rf_ram.memory[96][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__I0 (.I(\u_cpu.rf_ram.memory[96][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__A1 (.I(\u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__I2 (.I(\u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__A1 (.I(\u_cpu.rf_ram.memory[98][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__I2 (.I(\u_cpu.rf_ram.memory[98][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A1 (.I(\u_cpu.rf_ram.memory[98][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__I2 (.I(\u_cpu.rf_ram.memory[98][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__A1 (.I(\u_cpu.rf_ram.memory[98][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__I2 (.I(\u_cpu.rf_ram.memory[98][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__A1 (.I(\u_cpu.rf_ram.memory[98][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__I2 (.I(\u_cpu.rf_ram.memory[98][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A1 (.I(\u_cpu.rf_ram.memory[98][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__I2 (.I(\u_cpu.rf_ram.memory[98][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(\u_cpu.rf_ram.memory[99][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__I3 (.I(\u_cpu.rf_ram.memory[99][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A1 (.I(\u_cpu.rf_ram.memory[99][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__I3 (.I(\u_cpu.rf_ram.memory[99][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A1 (.I(\u_cpu.rf_ram.memory[99][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__I3 (.I(\u_cpu.rf_ram.memory[99][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A1 (.I(\u_cpu.rf_ram.memory[99][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__I3 (.I(\u_cpu.rf_ram.memory[99][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A1 (.I(\u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__I1 (.I(\u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__A1 (.I(\u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__I1 (.I(\u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__A1 (.I(\u_cpu.rf_ram.memory[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__I1 (.I(\u_cpu.rf_ram.memory[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A1 (.I(\u_cpu.rf_ram.memory[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__I1 (.I(\u_cpu.rf_ram.memory[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A1 (.I(\u_cpu.rf_ram.memory[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__I1 (.I(\u_cpu.rf_ram.memory[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A1 (.I(\u_cpu.rf_ram.memory[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__I1 (.I(\u_cpu.rf_ram.memory[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A1 (.I(\u_cpu.rf_ram.memory[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__I1 (.I(\u_cpu.rf_ram.memory[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A2 (.I(\u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__A2 (.I(\u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A2 (.I(\u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__D (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__A3 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A2 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__A2 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__A1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13039__I (.I(\u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout538_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout512_I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12057__CLK (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12056__CLK (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12052__CLK (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12055__CLK (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout8_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12777__CLK (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12773__CLK (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12772__CLK (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__CLK (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11832__CLK (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12778__CLK (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout12_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12776__CLK (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout11_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout13_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout9_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout10_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__CLK (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__CLK (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__CLK (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12058__CLK (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout15_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11799__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11795__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12779__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11828__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout18_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout19_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout16_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout17_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout20_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout14_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout21_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12060__CLK (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__CLK (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12038__CLK (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__CLK (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11948__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11947__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11956__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__CLK (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__CLK (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11952__CLK (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11951__CLK (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__CLK (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__CLK (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout25_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12036__CLK (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout24_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11972__CLK (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11971__CLK (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11965__CLK (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__CLK (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__CLK (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11968__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11967__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11966__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout28_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout29_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout30_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout27_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11802__CLK (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11812__CLK (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11801__CLK (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__CLK (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__CLK (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__CLK (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__CLK (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__CLK (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11811__CLK (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout34_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11954__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11938__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12793__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11970__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout38_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout32_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout22_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12141__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12135__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12023__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12022__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12014__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12021__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12015__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12013__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12006__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12005__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12683__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12682__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12681__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12680__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12672__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12671__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12430__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12429__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12426__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12132__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12151__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12142__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12134__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12493__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12150__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12148__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12140__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12011__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12003__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12072__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12071__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12070__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12068__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12133__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12025__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12017__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12012__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12085__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12084__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12083__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12073__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12024__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11936__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12074__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12010__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11944__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11943__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11935__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12792__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12789__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12090__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12026__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11942__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11923__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12790__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12139__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12131__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12152__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12145__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12166__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12155__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12169__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12163__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12156__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12154__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12146__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12138__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12164__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12168__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12160__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11777__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11776__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11900__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11895__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11894__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11887__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11886__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11774__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11771__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11849__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11856__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11841__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11840__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12820__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12804__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11847__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11846__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12781__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12780__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11861__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12805__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11864__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11851__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11836__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12841__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout114_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12842__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12839__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12826__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12823__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12783__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12737__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12733__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12732__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12725__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12724__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12731__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12730__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12828__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12819__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12812__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11810__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11809__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12728__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12727__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12726__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11806__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout126_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12831__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12830__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12829__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12708__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12693__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12715__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12714__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12713__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12709__CLK (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout134_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12834__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12770__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12769__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12768__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12766__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12751__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12750__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12649__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12648__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12647__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12639__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12752__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12638__CLK (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12636__CLK (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12646__CLK (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12619__CLK (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12618__CLK (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12736__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12735__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12734__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12620__CLK (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12712__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12711__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12710__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12634__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12613__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12645__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12635__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12617__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12614__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout156_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout153_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout154_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout157_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout151_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout152_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12652__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12630__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12628__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12616__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12615__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12654__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout159_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout158_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout160_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout150_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout161_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11641__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11639__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout164_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12791__CLK (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__CLK (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__CLK (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11789__CLK (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11869__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12595__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11882__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11792__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11790__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout167_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout168_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout163_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout165_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__CLK (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout170_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12765__CLK (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12764__CLK (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12593__CLK (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout173_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12594__CLK (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12592__CLK (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12591__CLK (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12590__CLK (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12915__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12911__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12917__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12667__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12660__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12507__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout175_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout176_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout177_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout172_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout174_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout178_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout171_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout179_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout169_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11875__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11880__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11879__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12553__CLK (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout183_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout181_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout182_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12179__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11881__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11874__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11873__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout184_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout187_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12552__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12551__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12510__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12509__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout190_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout186_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout188_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout191_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout185_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout192_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout180_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12688__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12657__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12633__CLK (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12902__CLK (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12651__CLK (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12650__CLK (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__CLK (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12914__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12913__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12912__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12307__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12306__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12305__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12304__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12303__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout198_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout199_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12907__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12903__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout200_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout196_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout197_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout201_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout194_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout195_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12906__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12904__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12653__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12629__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12627__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout204_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout205_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout202_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12759__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12302__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12762__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12761__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12758__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12760__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout207_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11629__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__CLK (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout209_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout210_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout208_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11636__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11922__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11915__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11733__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout213_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout214_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__CLK (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout212_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout215_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout211_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11730__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11729__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout217_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout218_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11918__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11921__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11920__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11916__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11984__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11979__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout220_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11988__CLK (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11987__CLK (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11994__CLK (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__CLK (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__CLK (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout223_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout224_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__CLK (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout222_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout226_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__CLK (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout219_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout227_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout216_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout228_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout206_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout229_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout193_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout230_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout162_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout231_I (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12433__CLK (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12432__CLK (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12431__CLK (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12425__CLK (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12424__CLK (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12434__CLK (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12421__CLK (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12420__CLK (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout233_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout234_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12659__CLK (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12435__CLK (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12473__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12492__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12491__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12490__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout237_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout238_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__CLK (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12479__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12494__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12480__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12478__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12484__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12488__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12487__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12486__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12485__CLK (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout242_I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout240_I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout241_I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout243_I (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout239_I (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout244_I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout235_I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout236_I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12417__CLK (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12416__CLK (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12413__CLK (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12441__CLK (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout246_I (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12444__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12415__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12414__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12442__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout249_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout250_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout247_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout248_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12458__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12462__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12456__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12459__CLK (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout253_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12545__CLK (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout252_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12544__CLK (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12512__CLK (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12297__CLK (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12272__CLK (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout254_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout255_I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout251_I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout256_I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout245_I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12100__CLK (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12191__CLK (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12190__CLK (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__CLK (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12187__CLK (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout260_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout261_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout258_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout259_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12624__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12621__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12622__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12463__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12116__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12115__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12103__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12101__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12099__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout264_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout265_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12625__CLK (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout263_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout266_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout262_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11780__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12194__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12193__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12192__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11786__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11890__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11897__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11896__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11889__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11888__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout270_I (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout271_I (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout268_I (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout269_I (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12106__CLK (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__CLK (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__CLK (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11781__CLK (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11779__CLK (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12121__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12120__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11785__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11910__CLK (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__CLK (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11908__CLK (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout273_I (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout274_I (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout275_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout276_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout272_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout277_I (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout267_I (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12957__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12945__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12472__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12958__CLK (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__CLK (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12236__CLK (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__CLK (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12944__CLK (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__CLK (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12232__CLK (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12231__CLK (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout281_I (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout282_I (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12119__CLK (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__CLK (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12943__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12234__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout287_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout288_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout285_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout286_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout289_I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout284_I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__CLK (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12110__CLK (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12109__CLK (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout291_I (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout292_I (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12204__CLK (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12203__CLK (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12196__CLK (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11706__CLK (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11704__CLK (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout295_I (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout296_I (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout293_I (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout294_I (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__CLK (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12198__CLK (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__CLK (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12205__CLK (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12197__CLK (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__CLK (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11763__CLK (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12218__CLK (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12210__CLK (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12202__CLK (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout300_I (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout301_I (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout298_I (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout299_I (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout302_I (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout297_I (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout303_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout290_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout304_I (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout278_I (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout305_I (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout257_I (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12513__CLK (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__CLK (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12516__CLK (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12515__CLK (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12514__CLK (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12560__CLK (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12559__CLK (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12565__CLK (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12564__CLK (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12563__CLK (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12562__CLK (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12561__CLK (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout310_I (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12522__CLK (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__CLK (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12519__CLK (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__CLK (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout309_I (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout311_I (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout307_I (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout308_I (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12555__CLK (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12279__CLK (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12278__CLK (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12556__CLK (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12554__CLK (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12296__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12275__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12274__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12935__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout313_I (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12495__CLK (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11734__CLK (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12299__CLK (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12276__CLK (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12273__CLK (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12542__CLK (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12541__CLK (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12540__CLK (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout316_I (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout317_I (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout318_I (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12587__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12586__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12585__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12277__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12946__CLK (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout319_I (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout314_I (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout315_I (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout320_I (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout312_I (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__CLK (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__CLK (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12524__CLK (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12523__CLK (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12521__CLK (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12531__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12530__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12529__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12528__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12527__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12575__CLK (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12574__CLK (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12573__CLK (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12532__CLK (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout324_I (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout325_I (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout322_I (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout323_I (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12584__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12581__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12571__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12578__CLK (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12577__CLK (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12576__CLK (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12533__CLK (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12580__CLK (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__CLK (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12535__CLK (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__CLK (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12579__CLK (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout329_I (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout330_I (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout327_I (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout328_I (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout331_I (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout326_I (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout332_I (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout321_I (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12857__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12956__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12948__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12856__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12852__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout336_I (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12094__CLK (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12092__CLK (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12091__CLK (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11736__CLK (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12096__CLK (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout337_I (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout334_I (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout335_I (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout340_I (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12952__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12951__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12950__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12949__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout339_I (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout341_I (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout338_I (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12097__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12217__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12216__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12199__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__CLK (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12222__CLK (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12098__CLK (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12225__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11767__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11766__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12253__CLK (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12249__CLK (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12248__CLK (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12221__CLK (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12219__CLK (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12256__CLK (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12255__CLK (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12254__CLK (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12220__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12345__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12344__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12341__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout350_I (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout351_I (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout348_I (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout349_I (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout352_I (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout347_I (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout353_I (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout342_I (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12266__CLK (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12264__CLK (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12260__CLK (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12259__CLK (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12258__CLK (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12244__CLK (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12243__CLK (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__CLK (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12269__CLK (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12265__CLK (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout359_I (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12263__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12262__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12261__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12257__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout361_I (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout362_I (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout358_I (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout360_I (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12335__CLK (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12334__CLK (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12353__CLK (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12352__CLK (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12351__CLK (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout366_I (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout363_I (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout367_I (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout357_I (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout368_I (.I(net369));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout354_I (.I(net369));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout369_I (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout333_I (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout370_I (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout306_I (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12182__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11899__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11898__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12181__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11914__CLK (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__CLK (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__CLK (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11724__CLK (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11723__CLK (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout375_I (.I(net377));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout376_I (.I(net377));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout372_I (.I(net377));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout373_I (.I(net377));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12932__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12931__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12930__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12934__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12929__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12933__CLK (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout378_I (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__CLK (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__CLK (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12293__CLK (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12289__CLK (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12288__CLK (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12281__CLK (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12280__CLK (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout380_I (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__CLK (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__CLK (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__CLK (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__CLK (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout382_I (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout383_I (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12925__CLK (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout381_I (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout384_I (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout379_I (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout385_I (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout377_I (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11702__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout390_I (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__CLK (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__CLK (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__CLK (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__CLK (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout389_I (.I(net392));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout391_I (.I(net392));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout387_I (.I(net392));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout388_I (.I(net392));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__CLK (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11755__CLK (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__CLK (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11762__CLK (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__CLK (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11650__CLK (.I(net395));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11649__CLK (.I(net395));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11648__CLK (.I(net395));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout393_I (.I(net395));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout394_I (.I(net395));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout395_I (.I(net397));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout396_I (.I(net397));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout392_I (.I(net397));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12283__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12282__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12291__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12290__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout399_I (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12295__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12294__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12287__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12285__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11661__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11647__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11657__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11716__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout403_I (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout404_I (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__CLK (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__CLK (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__CLK (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout405_I (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout401_I (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout402_I (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout406_I (.I(net407));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout398_I (.I(net407));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout400_I (.I(net407));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout407_I (.I(net408));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout397_I (.I(net408));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout408_I (.I(net409));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout386_I (.I(net409));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12798__CLK (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12797__CLK (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12796__CLK (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout410_I (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout411_I (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout414_I (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12803__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12802__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12801__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout416_I (.I(net418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout417_I (.I(net418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout412_I (.I(net418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout413_I (.I(net418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12034__CLK (.I(net419));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12033__CLK (.I(net419));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__CLK (.I(net419));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__CLK (.I(net419));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__CLK (.I(net419));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout419_I (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout420_I (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11983__CLK (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__CLK (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11981__CLK (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12369__CLK (.I(net422));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12368__CLK (.I(net422));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12367__CLK (.I(net422));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12366__CLK (.I(net422));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__CLK (.I(net422));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout424_I (.I(net426));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout425_I (.I(net426));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout422_I (.I(net426));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout423_I (.I(net426));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout426_I (.I(net427));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout421_I (.I(net427));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout427_I (.I(net428));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout418_I (.I(net428));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11744__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11743__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11751__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout429_I (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12895__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12894__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11747__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout432_I (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout433_I (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout430_I (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout431_I (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__CLK (.I(net435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12851__CLK (.I(net435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12848__CLK (.I(net435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12844__CLK (.I(net435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__CLK (.I(net435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12847__CLK (.I(net437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12901__CLK (.I(net437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12900__CLK (.I(net437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12899__CLK (.I(net437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__CLK (.I(net437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout437_I (.I(net439));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout438_I (.I(net439));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout435_I (.I(net439));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout436_I (.I(net439));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout439_I (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout434_I (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12598__CLK (.I(net441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12597__CLK (.I(net441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12360__CLK (.I(net441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12359__CLK (.I(net441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__CLK (.I(net441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12610__CLK (.I(net443));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12606__CLK (.I(net443));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12605__CLK (.I(net443));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout441_I (.I(net443));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout442_I (.I(net443));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12599__CLK (.I(net445));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__CLK (.I(net445));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__CLK (.I(net445));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__CLK (.I(net445));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__CLK (.I(net445));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12609__CLK (.I(net447));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__CLK (.I(net447));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__CLK (.I(net447));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout445_I (.I(net447));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout446_I (.I(net447));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout447_I (.I(net448));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout443_I (.I(net448));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout444_I (.I(net448));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout448_I (.I(net449));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout440_I (.I(net449));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout449_I (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout428_I (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout450_I (.I(net451));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout409_I (.I(net451));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__CLK (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__CLK (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12348__CLK (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12347__CLK (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11757__CLK (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout454_I (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12403__CLK (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12402__CLK (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12401__CLK (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12346__CLK (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11689__CLK (.I(net456));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__CLK (.I(net456));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12404__CLK (.I(net456));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11692__CLK (.I(net456));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11691__CLK (.I(net456));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout458_I (.I(net459));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12400__CLK (.I(net459));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout455_I (.I(net459));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout459_I (.I(net460));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout452_I (.I(net460));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout453_I (.I(net460));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__CLK (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout461_I (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__CLK (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__CLK (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout462_I (.I(net463));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11710__CLK (.I(net463));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__CLK (.I(net463));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__CLK (.I(net463));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12314__CLK (.I(net464));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__CLK (.I(net464));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11686__CLK (.I(net464));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__CLK (.I(net464));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__CLK (.I(net464));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12322__CLK (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__CLK (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12310__CLK (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__CLK (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout466_I (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12324__CLK (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout467_I (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout464_I (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout465_I (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout468_I (.I(net469));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout463_I (.I(net469));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout469_I (.I(net470));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout460_I (.I(net470));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12388__CLK (.I(net472));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12382__CLK (.I(net472));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12381__CLK (.I(net472));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12356__CLK (.I(net472));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12349__CLK (.I(net472));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12446__CLK (.I(net475));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12390__CLK (.I(net475));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12471__CLK (.I(net475));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout474_I (.I(net475));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout475_I (.I(net476));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout472_I (.I(net476));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout473_I (.I(net476));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12392__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12451__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12447__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12395__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12391__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout481_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout482_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout479_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout480_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout483_I (.I(net484));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout476_I (.I(net484));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12407__CLK (.I(net485));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12411__CLK (.I(net485));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12410__CLK (.I(net485));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12405__CLK (.I(net485));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12315__CLK (.I(net485));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12311__CLK (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12323__CLK (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12321__CLK (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12317__CLK (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__CLK (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout487_I (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout488_I (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout485_I (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout486_I (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12500__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12469__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12468__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12467__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12394__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12498__CLK (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12497__CLK (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12496__CLK (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout490_I (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout491_I (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12499__CLK (.I(net493));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout492_I (.I(net493));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout489_I (.I(net493));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout493_I (.I(net494));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout484_I (.I(net494));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout494_I (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout470_I (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12878__CLK (.I(net496));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12877__CLK (.I(net496));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12870__CLK (.I(net496));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__CLK (.I(net496));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12862__CLK (.I(net496));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12871__CLK (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12863__CLK (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__CLK (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout496_I (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout497_I (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12867__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12876__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12875__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12872__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12864__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12873__CLK (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12866__CLK (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12865__CLK (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12868__CLK (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout500_I (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12882__CLK (.I(net502));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12874__CLK (.I(net502));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout501_I (.I(net503));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout502_I (.I(net503));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout498_I (.I(net503));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout499_I (.I(net503));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__CLK (.I(net504));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout503_I (.I(net504));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout507_I (.I(net508));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout504_I (.I(net508));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout508_I (.I(net509));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout495_I (.I(net509));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout509_I (.I(net510));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout451_I (.I(net510));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout510_I (.I(net511));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout371_I (.I(net511));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout511_I (.I(net512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout232_I (.I(net512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12978__CLK (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12976__CLK (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12979__CLK (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout513_I (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12987__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12973__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12986__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12985__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12977__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12972__CLK (.I(net517));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12971__CLK (.I(net517));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12970__CLK (.I(net517));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12988__CLK (.I(net517));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout516_I (.I(net517));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12974__CLK (.I(net518));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout517_I (.I(net518));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout515_I (.I(net518));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12967__CLK (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12966__CLK (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12991__CLK (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12990__CLK (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12989__CLK (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12962__CLK (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12995__CLK (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12994__CLK (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12993__CLK (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12992__CLK (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout521_I (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout522_I (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout519_I (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout520_I (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout523_I (.I(net524));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout518_I (.I(net524));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12998__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13002__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13001__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12997__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12996__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13005__CLK (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13004__CLK (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13003__CLK (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout525_I (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout526_I (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13027__CLK (.I(net529));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12961__CLK (.I(net529));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12960__CLK (.I(net529));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout527_I (.I(net529));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout528_I (.I(net529));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13010__CLK (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13009__CLK (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13008__CLK (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13013__CLK (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13012__CLK (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13017__CLK (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13016__CLK (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13015__CLK (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout530_I (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout531_I (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13029__CLK (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__CLKN (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13022__CLK (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13021__CLK (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13020__CLK (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout534_I (.I(net535));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13026__CLK (.I(net535));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13025__CLK (.I(net535));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13024__CLK (.I(net535));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13023__CLK (.I(net535));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13038__I (.I(net536));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout535_I (.I(net536));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout532_I (.I(net536));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout533_I (.I(net536));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout536_I (.I(net537));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13028__CLK (.I(net537));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout529_I (.I(net537));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout537_I (.I(net538));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout524_I (.I(net538));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1758 ();
 assign io_oeb[0] = net539;
 assign io_oeb[1] = net540;
 assign io_oeb[2] = net541;
 assign io_oeb[3] = net542;
 assign io_oeb[4] = net543;
 assign io_out[2] = net544;
 assign io_out[3] = net545;
 assign io_out[4] = net546;
endmodule

